// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 15 2024 15:29:08

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "State_Machine_Project_Top" view "INTERFACE"

module State_Machine_Project_Top (
    o_Segment2_D,
    o_LED_3,
    i_Switch_4,
    i_Clk,
    o_Segment2_G,
    o_Segment2_C,
    o_LED_2,
    i_Switch_1,
    o_Segment2_F,
    o_Segment2_B,
    o_LED_1,
    i_Switch_2,
    o_Segment2_E,
    o_Segment2_A,
    o_LED_4,
    i_Switch_3);

    output o_Segment2_D;
    output o_LED_3;
    input i_Switch_4;
    input i_Clk;
    output o_Segment2_G;
    output o_Segment2_C;
    output o_LED_2;
    input i_Switch_1;
    output o_Segment2_F;
    output o_Segment2_B;
    output o_LED_1;
    input i_Switch_2;
    output o_Segment2_E;
    output o_Segment2_A;
    output o_LED_4;
    input i_Switch_3;

    wire N__8739;
    wire N__8738;
    wire N__8737;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8719;
    wire N__8718;
    wire N__8717;
    wire N__8710;
    wire N__8709;
    wire N__8708;
    wire N__8701;
    wire N__8700;
    wire N__8699;
    wire N__8692;
    wire N__8691;
    wire N__8690;
    wire N__8683;
    wire N__8682;
    wire N__8681;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8665;
    wire N__8664;
    wire N__8663;
    wire N__8656;
    wire N__8655;
    wire N__8654;
    wire N__8647;
    wire N__8646;
    wire N__8645;
    wire N__8638;
    wire N__8637;
    wire N__8636;
    wire N__8629;
    wire N__8628;
    wire N__8627;
    wire N__8620;
    wire N__8619;
    wire N__8618;
    wire N__8611;
    wire N__8610;
    wire N__8609;
    wire N__8602;
    wire N__8601;
    wire N__8600;
    wire N__8583;
    wire N__8582;
    wire N__8579;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8540;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8530;
    wire N__8523;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8489;
    wire N__8486;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8478;
    wire N__8477;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8451;
    wire N__8450;
    wire N__8449;
    wire N__8448;
    wire N__8447;
    wire N__8446;
    wire N__8445;
    wire N__8444;
    wire N__8443;
    wire N__8442;
    wire N__8441;
    wire N__8440;
    wire N__8439;
    wire N__8438;
    wire N__8437;
    wire N__8436;
    wire N__8435;
    wire N__8434;
    wire N__8433;
    wire N__8432;
    wire N__8431;
    wire N__8430;
    wire N__8429;
    wire N__8428;
    wire N__8427;
    wire N__8426;
    wire N__8425;
    wire N__8424;
    wire N__8423;
    wire N__8422;
    wire N__8421;
    wire N__8420;
    wire N__8419;
    wire N__8418;
    wire N__8417;
    wire N__8416;
    wire N__8415;
    wire N__8414;
    wire N__8413;
    wire N__8412;
    wire N__8411;
    wire N__8410;
    wire N__8409;
    wire N__8408;
    wire N__8407;
    wire N__8406;
    wire N__8405;
    wire N__8404;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8300;
    wire N__8299;
    wire N__8296;
    wire N__8291;
    wire N__8286;
    wire N__8285;
    wire N__8282;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8265;
    wire N__8264;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8252;
    wire N__8247;
    wire N__8246;
    wire N__8245;
    wire N__8242;
    wire N__8237;
    wire N__8232;
    wire N__8231;
    wire N__8230;
    wire N__8227;
    wire N__8222;
    wire N__8217;
    wire N__8214;
    wire N__8213;
    wire N__8212;
    wire N__8209;
    wire N__8204;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8174;
    wire N__8171;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8154;
    wire N__8153;
    wire N__8152;
    wire N__8151;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8133;
    wire N__8132;
    wire N__8131;
    wire N__8130;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8088;
    wire N__8085;
    wire N__8084;
    wire N__8083;
    wire N__8080;
    wire N__8075;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8063;
    wire N__8062;
    wire N__8059;
    wire N__8054;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8031;
    wire N__8028;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8013;
    wire N__8010;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7995;
    wire N__7992;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7949;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7920;
    wire N__7917;
    wire N__7916;
    wire N__7915;
    wire N__7908;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7884;
    wire N__7883;
    wire N__7882;
    wire N__7875;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7857;
    wire N__7856;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7827;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7815;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7803;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7791;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7779;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7767;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7755;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7724;
    wire N__7719;
    wire N__7716;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7698;
    wire N__7695;
    wire N__7694;
    wire N__7693;
    wire N__7690;
    wire N__7689;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7671;
    wire N__7668;
    wire N__7667;
    wire N__7664;
    wire N__7663;
    wire N__7660;
    wire N__7657;
    wire N__7654;
    wire N__7647;
    wire N__7646;
    wire N__7645;
    wire N__7644;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7628;
    wire N__7627;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7605;
    wire N__7604;
    wire N__7603;
    wire N__7602;
    wire N__7601;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7583;
    wire N__7582;
    wire N__7581;
    wire N__7578;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7567;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7556;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7528;
    wire N__7523;
    wire N__7520;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7490;
    wire N__7489;
    wire N__7486;
    wire N__7481;
    wire N__7478;
    wire N__7477;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7366;
    wire N__7359;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7332;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7310;
    wire N__7309;
    wire N__7306;
    wire N__7301;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7289;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7279;
    wire N__7274;
    wire N__7269;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7257;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7242;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7230;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7202;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7185;
    wire N__7182;
    wire N__7181;
    wire N__7180;
    wire N__7177;
    wire N__7172;
    wire N__7167;
    wire N__7164;
    wire N__7163;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7146;
    wire N__7143;
    wire N__7142;
    wire N__7141;
    wire N__7138;
    wire N__7133;
    wire N__7128;
    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7104;
    wire N__7101;
    wire N__7100;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7083;
    wire N__7080;
    wire N__7079;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7056;
    wire N__7053;
    wire N__7052;
    wire N__7051;
    wire N__7048;
    wire N__7043;
    wire N__7038;
    wire N__7035;
    wire N__7034;
    wire N__7033;
    wire N__7030;
    wire N__7025;
    wire N__7020;
    wire N__7019;
    wire N__7018;
    wire N__7015;
    wire N__7010;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6996;
    wire N__6995;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6983;
    wire N__6980;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6963;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6951;
    wire N__6948;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6933;
    wire N__6930;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6918;
    wire N__6915;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6903;
    wire N__6900;
    wire N__6899;
    wire N__6896;
    wire N__6895;
    wire N__6892;
    wire N__6887;
    wire N__6882;
    wire N__6879;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6857;
    wire N__6856;
    wire N__6853;
    wire N__6848;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6816;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6771;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6725;
    wire N__6724;
    wire N__6721;
    wire N__6716;
    wire N__6711;
    wire N__6710;
    wire N__6709;
    wire N__6706;
    wire N__6701;
    wire N__6696;
    wire N__6695;
    wire N__6694;
    wire N__6691;
    wire N__6686;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6671;
    wire N__6670;
    wire N__6667;
    wire N__6664;
    wire N__6659;
    wire N__6654;
    wire N__6653;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6636;
    wire N__6635;
    wire N__6632;
    wire N__6631;
    wire N__6628;
    wire N__6623;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6594;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6582;
    wire N__6579;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6571;
    wire N__6570;
    wire N__6569;
    wire N__6568;
    wire N__6567;
    wire N__6566;
    wire N__6565;
    wire N__6564;
    wire N__6563;
    wire N__6562;
    wire N__6557;
    wire N__6554;
    wire N__6549;
    wire N__6542;
    wire N__6537;
    wire N__6532;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6492;
    wire N__6491;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6465;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6450;
    wire N__6449;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6432;
    wire N__6429;
    wire N__6428;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6411;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6315;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6291;
    wire N__6288;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6173;
    wire N__6172;
    wire N__6169;
    wire N__6164;
    wire N__6163;
    wire N__6162;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6147;
    wire N__6138;
    wire N__6135;
    wire N__6134;
    wire N__6133;
    wire N__6128;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6114;
    wire N__6113;
    wire N__6112;
    wire N__6109;
    wire N__6108;
    wire N__6107;
    wire N__6104;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6090;
    wire N__6089;
    wire N__6088;
    wire N__6087;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6070;
    wire N__6067;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6040;
    wire N__6027;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6002;
    wire N__6001;
    wire N__6000;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5985;
    wire N__5976;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5961;
    wire N__5960;
    wire N__5959;
    wire N__5958;
    wire N__5957;
    wire N__5956;
    wire N__5953;
    wire N__5948;
    wire N__5941;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5921;
    wire N__5916;
    wire N__5915;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5898;
    wire N__5895;
    wire N__5894;
    wire N__5889;
    wire N__5886;
    wire N__5885;
    wire N__5884;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5876;
    wire N__5873;
    wire N__5872;
    wire N__5871;
    wire N__5870;
    wire N__5869;
    wire N__5868;
    wire N__5867;
    wire N__5866;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5854;
    wire N__5851;
    wire N__5846;
    wire N__5843;
    wire N__5838;
    wire N__5835;
    wire N__5834;
    wire N__5829;
    wire N__5826;
    wire N__5817;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5793;
    wire N__5790;
    wire N__5789;
    wire N__5788;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5772;
    wire N__5769;
    wire N__5768;
    wire N__5767;
    wire N__5766;
    wire N__5765;
    wire N__5764;
    wire N__5759;
    wire N__5756;
    wire N__5751;
    wire N__5750;
    wire N__5749;
    wire N__5748;
    wire N__5747;
    wire N__5746;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5719;
    wire N__5706;
    wire N__5703;
    wire N__5702;
    wire N__5701;
    wire N__5698;
    wire N__5693;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5681;
    wire N__5678;
    wire N__5677;
    wire N__5676;
    wire N__5673;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5663;
    wire N__5662;
    wire N__5661;
    wire N__5660;
    wire N__5659;
    wire N__5658;
    wire N__5657;
    wire N__5656;
    wire N__5655;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5643;
    wire N__5638;
    wire N__5635;
    wire N__5628;
    wire N__5619;
    wire N__5604;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5585;
    wire N__5584;
    wire N__5581;
    wire N__5576;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5546;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5531;
    wire N__5530;
    wire N__5529;
    wire N__5526;
    wire N__5521;
    wire N__5516;
    wire N__5511;
    wire N__5510;
    wire N__5509;
    wire N__5508;
    wire N__5505;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5493;
    wire N__5490;
    wire N__5481;
    wire N__5480;
    wire N__5475;
    wire N__5474;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5457;
    wire N__5456;
    wire N__5455;
    wire N__5454;
    wire N__5453;
    wire N__5452;
    wire N__5443;
    wire N__5440;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5426;
    wire N__5425;
    wire N__5424;
    wire N__5421;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5394;
    wire N__5393;
    wire N__5392;
    wire N__5391;
    wire N__5390;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5379;
    wire N__5376;
    wire N__5373;
    wire N__5372;
    wire N__5363;
    wire N__5360;
    wire N__5355;
    wire N__5354;
    wire N__5351;
    wire N__5350;
    wire N__5347;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5322;
    wire N__5321;
    wire N__5320;
    wire N__5319;
    wire N__5318;
    wire N__5317;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5288;
    wire N__5287;
    wire N__5286;
    wire N__5283;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5260;
    wire N__5257;
    wire N__5250;
    wire N__5247;
    wire N__5246;
    wire N__5245;
    wire N__5244;
    wire N__5243;
    wire N__5242;
    wire N__5241;
    wire N__5238;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5222;
    wire N__5221;
    wire N__5220;
    wire N__5217;
    wire N__5212;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5173;
    wire N__5170;
    wire N__5169;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5157;
    wire N__5148;
    wire N__5147;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5127;
    wire N__5126;
    wire N__5125;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5106;
    wire N__5103;
    wire N__5100;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5046;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5031;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5009;
    wire N__5008;
    wire N__5001;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4976;
    wire N__4975;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4925;
    wire N__4924;
    wire N__4923;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4909;
    wire N__4902;
    wire N__4901;
    wire N__4900;
    wire N__4897;
    wire N__4892;
    wire N__4887;
    wire N__4886;
    wire N__4885;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4836;
    wire N__4833;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4818;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4776;
    wire N__4773;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4761;
    wire N__4758;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4746;
    wire N__4743;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4731;
    wire N__4728;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4713;
    wire N__4710;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4698;
    wire N__4695;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4680;
    wire N__4677;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4665;
    wire N__4662;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4647;
    wire N__4644;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4632;
    wire N__4629;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4617;
    wire N__4614;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4599;
    wire N__4596;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4581;
    wire N__4578;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4566;
    wire N__4563;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4551;
    wire N__4548;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4536;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4509;
    wire N__4506;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4476;
    wire N__4473;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4440;
    wire N__4437;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4410;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4370;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4358;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4280;
    wire N__4279;
    wire N__4276;
    wire N__4275;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4254;
    wire N__4253;
    wire N__4252;
    wire N__4251;
    wire N__4250;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4232;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4209;
    wire N__4208;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4195;
    wire N__4192;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4175;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4158;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4127;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4104;
    wire N__4103;
    wire N__4100;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4076;
    wire N__4075;
    wire N__4072;
    wire N__4067;
    wire N__4062;
    wire N__4061;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4023;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4011;
    wire N__4010;
    wire N__4009;
    wire N__4006;
    wire N__4001;
    wire N__3996;
    wire N__3995;
    wire N__3990;
    wire N__3987;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3951;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3923;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3900;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3888;
    wire N__3885;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3870;
    wire N__3867;
    wire N__3866;
    wire N__3865;
    wire N__3862;
    wire N__3857;
    wire N__3852;
    wire N__3849;
    wire N__3846;
    wire N__3845;
    wire N__3844;
    wire N__3841;
    wire N__3836;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire GNDG0;
    wire VCCG0;
    wire \Debounce_SW1.r_Count12_i ;
    wire \Debounce_SW1.N_28_1_cascade_ ;
    wire \Debounce_SW1.N_28_1 ;
    wire \Debounce_SW1.N_28 ;
    wire \Debounce_SW1.un1_r_Count_8lto17_i_3 ;
    wire \Debounce_SW1.r_Count13_10_cascade_ ;
    wire \Debounce_SW1.N_30 ;
    wire \Debounce_SW1.r_CountZ0Z_1 ;
    wire bfn_1_11_0_;
    wire \Debounce_SW1.r_CountZ0Z_2 ;
    wire \Debounce_SW1.r_Count_1_cry_1 ;
    wire \Debounce_SW1.r_CountZ0Z_3 ;
    wire \Debounce_SW1.r_Count_1_cry_2 ;
    wire \Debounce_SW1.r_CountZ0Z_4 ;
    wire \Debounce_SW1.r_Count_1_cry_3 ;
    wire \Debounce_SW1.r_Count_1_cry_4 ;
    wire \Debounce_SW1.r_CountZ0Z_6 ;
    wire \Debounce_SW1.r_Count_1_cry_5 ;
    wire \Debounce_SW1.r_Count_1_cry_6 ;
    wire \Debounce_SW1.r_CountZ0Z_8 ;
    wire \Debounce_SW1.r_Count_1_cry_7 ;
    wire \Debounce_SW1.r_Count_1_cry_8 ;
    wire bfn_1_12_0_;
    wire \Debounce_SW1.r_Count_1_cry_9 ;
    wire \Debounce_SW1.r_CountZ0Z_11 ;
    wire \Debounce_SW1.r_Count_1_cry_10 ;
    wire \Debounce_SW1.r_Count_1_cry_11 ;
    wire \Debounce_SW1.r_Count_1_cry_12 ;
    wire \Debounce_SW1.r_Count_1_cry_13 ;
    wire \Debounce_SW1.r_Count_1_cry_14 ;
    wire \Debounce_SW1.r_Count_1_cry_15 ;
    wire \Debounce_SW1.r_Count_1_cry_16 ;
    wire bfn_1_13_0_;
    wire \Debounce_SW1.r_CountZ0Z_0 ;
    wire \Debounce_SW1.r_Count12_i_g ;
    wire \Debounce_SW1.r_CountZ0Z_17 ;
    wire \Debounce_SW1.r_CountZ0Z_7 ;
    wire \Debounce_SW1.r_Count13_10 ;
    wire \Debounce_SW1.r_Count13_0_a7_4_cascade_ ;
    wire \Debounce_SW1.r_CountZ0Z_5 ;
    wire i_Switch_1_c;
    wire \Debounce_SW1.r_Count13_0_a7_7 ;
    wire \Debounce_SW1.r_Count13_0_a7_8_cascade_ ;
    wire \Debounce_SW1.r_CountZ0Z_16 ;
    wire \Debounce_SW1.r_CountZ0Z_12 ;
    wire \Debounce_SW1.un1_r_Count_8lto17_i_2 ;
    wire \Debounce_SW1.r_CountZ0Z_15 ;
    wire \Debounce_SW1.r_CountZ0Z_14 ;
    wire \Debounce_SW1.r_Count13_0_a7_0 ;
    wire \Debounce_SW1.r_CountZ0Z_10 ;
    wire \Debounce_SW1.r_CountZ0Z_9 ;
    wire \Debounce_SW1.r_CountZ0Z_13 ;
    wire \Debounce_SW1.N_28_2 ;
    wire \Game_Inst.Count_Inst.o_Toggle3_14 ;
    wire \Game_Inst.Count_Inst.o_Toggle3_13_cascade_ ;
    wire \Game_Inst.Count_Inst.o_Toggle3_12 ;
    wire \Game_Inst.Count_Inst.o_Toggle3_15 ;
    wire \Game_Inst.N_334_0_cascade_ ;
    wire \Game_Inst.N_249_0_cascade_ ;
    wire \Game_Inst.Count_Inst.r_Counter_RNIGDO97Z0Z_16 ;
    wire \Game_Inst.Count_Inst.o_Toggle3_17 ;
    wire \Game_Inst.Count_Inst.o_Toggle3_21 ;
    wire \Game_Inst.Count_Inst.o_Toggle3_17_cascade_ ;
    wire \Game_Inst.Count_Inst.o_Toggle3_16 ;
    wire \Game_Inst.N_249_0 ;
    wire \Game_Inst.Count_Inst.o_Toggle3_cascade_ ;
    wire \Game_Inst.r_SM_Main_ns_i_0_0_cascade_ ;
    wire \Game_Inst.r_SM_Main_ns_i_1_0_cascade_ ;
    wire \Game_Inst.r_SM_Main_ns_i_2_0_cascade_ ;
    wire \Game_Inst.N_338 ;
    wire \Game_Inst.r_SM_Main_ns_i_m2_ns_1_0 ;
    wire \Game_Inst.N_260_0_cascade_ ;
    wire \Game_Inst.N_260_0 ;
    wire r_Hex_Encoding_i_1;
    wire r_Hex_Encoding_i_5;
    wire r_Hex_Encoding_i_6;
    wire r_Hex_Encoding_i_3;
    wire r_Hex_Encoding_i_0;
    wire r_Hex_Encoding_i_4;
    wire bfn_5_4_0_;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_2 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_1 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_3 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_2 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_4 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_3 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_5 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_4 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_6 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_5 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_7 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_6 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_8 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_7 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_8 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_9 ;
    wire bfn_5_5_0_;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_10 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_9 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_11 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_10 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_12 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_11 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_13 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_12 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_14 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_13 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_15 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_14 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_16 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_15 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_16 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_17 ;
    wire bfn_5_6_0_;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_18 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_17 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_19 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_18 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_20 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_19 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_21 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_20 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_22 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_21 ;
    wire \Game_Inst.Count_Inst.un3_r_Counter_cry_22 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_23 ;
    wire \Game_Inst.r_SM_Main_ns_i_a4_0_0 ;
    wire \Game_Inst.r_SM_Main_ns_i_0_1_cascade_ ;
    wire \Game_Inst.r_SM_Main_ns_i_2_1_cascade_ ;
    wire \Game_Inst.r_SM_Main_ns_i_a4_0_1_1 ;
    wire \Game_Inst.w_Toggle ;
    wire \Game_Inst.r_ToggleZ0 ;
    wire \Game_Inst.r_SM_Main7 ;
    wire \Game_Inst.r_SM_Main_0_sqmuxa_2_1_cascade_ ;
    wire \Game_Inst.N_345 ;
    wire \Game_Inst.N_345_cascade_ ;
    wire \Game_Inst.SUM_i_0_1_cascade_ ;
    wire \Game_Inst.N_333_0 ;
    wire \Game_Inst.r_Index16_NE_1_cascade_ ;
    wire \Game_Inst.N_330_li ;
    wire \Game_Inst.N_330_li_cascade_ ;
    wire \Game_Inst.r_SM_Main_0_sqmuxa_1 ;
    wire \Game_Inst.r_Button_DVZ0 ;
    wire \Game_Inst.r_SM_Main_98_d_cascade_ ;
    wire \Game_Inst.o_Score_RNO_0Z0Z_0 ;
    wire bfn_5_10_0_;
    wire \Game_Inst.un1_o_Score_cry_0 ;
    wire \Game_Inst.o_Score_RNO_0Z0Z_2 ;
    wire \Game_Inst.un1_o_Score_cry_1 ;
    wire \Game_Inst.un1_o_Score_cry_2 ;
    wire \Game_Inst.o_Score_RNO_0Z0Z_3_cascade_ ;
    wire \Game_Inst.N_287_0_cascade_ ;
    wire \Game_Inst.N_262_0 ;
    wire \Game_Inst.o_Score_RNO_0Z0Z_1 ;
    wire \Game_Inst.N_287_0 ;
    wire \Game_Inst.o_Score_0_sqmuxa ;
    wire \Game_Inst.N_310 ;
    wire w_Score_1;
    wire w_Score_2;
    wire w_Score_3;
    wire w_Score_0;
    wire r_Hex_Encoding_i_2;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_0 ;
    wire \Game_Inst.Count_Inst.r_CounterZ0Z_1 ;
    wire \Game_Inst.Count_Inst.N_213_g ;
    wire \Game_Inst.r_SM_Main_100_d_cascade_ ;
    wire Game_Inst_o_LED_1_0_i;
    wire \Game_Inst.N_334_0 ;
    wire \Game_Inst.r_SM_Main_0_sqmuxa_2_1 ;
    wire \Game_Inst.N_335_0 ;
    wire \Game_Inst.r_SM_Main_ns_i_0_2 ;
    wire \Game_Inst.r_SM_MainZ0Z_0 ;
    wire \Game_Inst.N_275_0 ;
    wire \Game_Inst.N_275_0_cascade_ ;
    wire \Game_Inst.N_268_0_cascade_ ;
    wire \Game_Inst.r_Index_0_sqmuxa ;
    wire \Game_Inst.r_Pattern_1__RNIB13IZ0Z_0_cascade_ ;
    wire \Game_Inst.r_Pattern_2__RNIFHRIZ0Z_0 ;
    wire \Game_Inst.SUM_i_o3_1_0 ;
    wire \Game_Inst.un1_r_Pattern_0__7_ns_1_0 ;
    wire \Game_Inst.r_IndexZ1Z_1 ;
    wire \Game_Inst.N_276_0 ;
    wire \Game_Inst.r_IndexZ0Z_2 ;
    wire \Game_Inst.r_Pattern_5__RNIL3KJZ0Z_1_cascade_ ;
    wire \Game_Inst.un1_r_Pattern_0__7_ns_1_1 ;
    wire \Game_Inst.N_31_cascade_ ;
    wire \Game_Inst.un1_r_Pattern_0__1_i_0 ;
    wire \Game_Inst.N_311 ;
    wire \Game_Inst.r_SM_MainZ0Z_2 ;
    wire \Game_Inst.un1_r_Pattern_0__1_i_0_cascade_ ;
    wire \Game_Inst.N_309 ;
    wire \Game_Inst.r_SM_MainZ0Z_1 ;
    wire \Game_Inst.N_269_0_cascade_ ;
    wire \Game_Inst.N_314 ;
    wire \Game_Inst.r_SwitchZ0Z_4 ;
    wire \Game_Inst.r_Button_IDZ0Z_0 ;
    wire \Game_Inst.N_270_li ;
    wire \Game_Inst.r_SwitchZ0Z_1 ;
    wire w_Switch_1;
    wire \Game_Inst.r_Button_IDZ0Z_1 ;
    wire bfn_6_13_0_;
    wire \Debounce_SW2.r_Count_1_cry_1 ;
    wire \Debounce_SW2.r_Count_1_cry_2 ;
    wire \Debounce_SW2.r_Count_1_cry_3 ;
    wire \Debounce_SW2.r_Count_1_cry_4 ;
    wire \Debounce_SW2.r_Count_1_cry_5 ;
    wire \Debounce_SW2.r_Count_1_cry_6 ;
    wire \Debounce_SW2.r_Count_1_cry_7 ;
    wire \Debounce_SW2.r_Count_1_cry_8 ;
    wire bfn_6_14_0_;
    wire \Debounce_SW2.r_Count_1_cry_9 ;
    wire \Debounce_SW2.r_Count_1_cry_10 ;
    wire \Debounce_SW2.r_Count_1_cry_11 ;
    wire \Debounce_SW2.r_Count_1_cry_12 ;
    wire \Debounce_SW2.r_Count_1_cry_13 ;
    wire \Debounce_SW2.r_Count_1_cry_14 ;
    wire \Debounce_SW2.r_Count_1_cry_15 ;
    wire \Debounce_SW2.r_Count_1_cry_16 ;
    wire bfn_6_15_0_;
    wire \Debounce_SW4.r_Count12_i ;
    wire i_Switch_4_c;
    wire \Debounce_SW4.r_Count13_10_2 ;
    wire \Debounce_SW4.r_Count13_9_cascade_ ;
    wire \Debounce_SW4.r_Count13_1 ;
    wire \Debounce_SW4.r_Count13_1_cascade_ ;
    wire \Debounce_SW4.un1_r_Count_8lt11_0_cascade_ ;
    wire \Debounce_SW4.un1_r_Count_8lt17 ;
    wire \Debounce_SW4.un1_r_Count_8lto11_1 ;
    wire \Debounce_SW4.un1_r_Count_8lto17_2 ;
    wire \Debounce_SW4.r_Count13_5 ;
    wire \Debounce_SW4.r_Count13_6 ;
    wire \Game_Inst.r_Pattern_1__RNID33IZ0Z_1 ;
    wire \Game_Inst.r_Pattern_2__RNIHJRIZ0Z_1 ;
    wire \Game_Inst.r_Pattern_0_Z0Z_1 ;
    wire \Game_Inst.r_Pattern_2_Z0Z_1 ;
    wire \Game_Inst.r_Pattern_3_Z0Z_1 ;
    wire \Game_Inst.r_Pattern_1_Z0Z_1 ;
    wire \Game_Inst.r_Pattern_0_Z0Z_0 ;
    wire \Game_Inst.r_Pattern_1_Z0Z_0 ;
    wire \Game_Inst.r_Pattern_2_Z0Z_0 ;
    wire \Game_Inst.r_Pattern_3_Z0Z_0 ;
    wire \Game_Inst.w_LFSR_Data_3 ;
    wire \Game_Inst.r_Pattern_6__RNIPJCKZ0Z_1 ;
    wire \Game_Inst.w_LFSR_Data_4 ;
    wire \Game_Inst.r_Pattern_6__RNINHCKZ0Z_0 ;
    wire \Game_Inst.w_LFSR_Data_1 ;
    wire \Game_Inst.w_LFSR_Data_2 ;
    wire \Game_Inst.r_IndexZ0Z_0 ;
    wire \Game_Inst.r_Pattern_5__RNIJ1KJZ0Z_0 ;
    wire \Game_Inst.un1_i_Switch_4_1 ;
    wire \Game_Inst.r_Button_ID_2_0 ;
    wire \Debounce_SW2.r_Count13_0_a7_7 ;
    wire \Debounce_SW2.r_CountZ0Z_2 ;
    wire \Debounce_SW2.r_CountZ0Z_3 ;
    wire \Debounce_SW2.r_CountZ0Z_6 ;
    wire \Debounce_SW2.r_Count13_10_cascade_ ;
    wire \Debounce_SW2.r_CountZ0Z_4 ;
    wire \Debounce_SW2.r_CountZ0Z_11 ;
    wire \Debounce_SW2.r_CountZ0Z_8 ;
    wire \Debounce_SW2.r_Count13_10 ;
    wire \Debounce_SW2.r_CountZ0Z_5 ;
    wire \Debounce_SW2.r_Count13_0_a7_8 ;
    wire \Debounce_SW2.r_Count13_0_a7_0 ;
    wire \Debounce_SW2.r_CountZ0Z_9 ;
    wire \Debounce_SW2.r_CountZ0Z_10 ;
    wire \Debounce_SW2.N_23_2 ;
    wire \Debounce_SW2.N_23_1 ;
    wire \Debounce_SW2.N_23_2_cascade_ ;
    wire \Debounce_SW2.N_25 ;
    wire i_Switch_2_c;
    wire \Debounce_SW2.N_23_cascade_ ;
    wire \Debounce_SW2.r_Count12_i ;
    wire \Debounce_SW2.r_CountZ0Z_15 ;
    wire \Debounce_SW2.r_CountZ0Z_13 ;
    wire \Debounce_SW2.r_CountZ0Z_14 ;
    wire \Debounce_SW2.un1_r_Count_8lto17_i_2_cascade_ ;
    wire \Debounce_SW2.un1_r_Count_8lto17_i_3 ;
    wire \Debounce_SW2.r_CountZ0Z_16 ;
    wire \Debounce_SW2.r_CountZ0Z_17 ;
    wire \Debounce_SW2.r_CountZ0Z_7 ;
    wire \Debounce_SW2.r_CountZ0Z_12 ;
    wire \Debounce_SW2.r_Count13_0_a7_4 ;
    wire \Debounce_SW4.r_Count13_10 ;
    wire \Debounce_SW4.r_CountZ0Z_1 ;
    wire bfn_8_5_0_;
    wire \Debounce_SW4.r_CountZ0Z_2 ;
    wire \Debounce_SW4.r_Count_1_cry_1 ;
    wire \Debounce_SW4.r_CountZ0Z_3 ;
    wire \Debounce_SW4.r_Count_1_cry_2 ;
    wire \Debounce_SW4.r_CountZ0Z_4 ;
    wire \Debounce_SW4.r_Count_1_cry_3 ;
    wire \Debounce_SW4.r_CountZ0Z_5 ;
    wire \Debounce_SW4.r_Count_1_cry_4 ;
    wire \Debounce_SW4.r_CountZ0Z_6 ;
    wire \Debounce_SW4.r_Count_1_cry_5 ;
    wire \Debounce_SW4.r_CountZ0Z_7 ;
    wire \Debounce_SW4.r_Count_1_cry_6 ;
    wire \Debounce_SW4.r_CountZ0Z_8 ;
    wire \Debounce_SW4.r_Count_1_cry_7 ;
    wire \Debounce_SW4.r_Count_1_cry_8 ;
    wire \Debounce_SW4.r_CountZ0Z_9 ;
    wire bfn_8_6_0_;
    wire \Debounce_SW4.r_CountZ0Z_10 ;
    wire \Debounce_SW4.r_Count_1_cry_9 ;
    wire \Debounce_SW4.r_CountZ0Z_11 ;
    wire \Debounce_SW4.r_Count_1_cry_10 ;
    wire \Debounce_SW4.r_CountZ0Z_12 ;
    wire \Debounce_SW4.r_Count_1_cry_11 ;
    wire \Debounce_SW4.r_CountZ0Z_13 ;
    wire \Debounce_SW4.r_Count_1_cry_12 ;
    wire \Debounce_SW4.r_CountZ0Z_14 ;
    wire \Debounce_SW4.r_Count_1_cry_13 ;
    wire \Debounce_SW4.r_CountZ0Z_15 ;
    wire \Debounce_SW4.r_Count_1_cry_14 ;
    wire \Debounce_SW4.r_CountZ0Z_16 ;
    wire \Debounce_SW4.r_Count_1_cry_15 ;
    wire \Debounce_SW4.r_Count_1_cry_16 ;
    wire bfn_8_7_0_;
    wire \Debounce_SW4.r_CountZ0Z_17 ;
    wire \Game_Inst.w_LFSR_Data_7 ;
    wire \Game_Inst.w_LFSR_Data_5 ;
    wire \Game_Inst.w_LFSR_Data_6 ;
    wire \Game_Inst.w_LFSR_Data_8 ;
    wire \Game_Inst.r_Pattern_4_Z0Z_0 ;
    wire \Game_Inst.r_Pattern_4_Z0Z_1 ;
    wire \Game_Inst.r_Pattern_5_Z0Z_0 ;
    wire \Game_Inst.r_Pattern_5_Z0Z_1 ;
    wire \Game_Inst.r_Pattern_6_Z0Z_0 ;
    wire \Game_Inst.r_Pattern_6_Z0Z_1 ;
    wire \Game_Inst.r_Pattern_7_Z0Z_0 ;
    wire \Game_Inst.r_Pattern_7_Z0Z_1 ;
    wire \Game_Inst.r_SM_Main_98_d ;
    wire \Game_Inst.r_Button_ID_2_sm0_0 ;
    wire \Game_Inst.r_SwitchZ0Z_2 ;
    wire \Game_Inst.r_SwitchZ0Z_3 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_19 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_21 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_20 ;
    wire \Game_Inst.w_LFSR_Data_0 ;
    wire \Debounce_SW2.r_CountZ0Z_0 ;
    wire \Debounce_SW2.r_CountZ0Z_1 ;
    wire \Debounce_SW2.r_Count12_i_g ;
    wire \Debounce_SW4.r_CountZ0Z_0 ;
    wire \Debounce_SW4.r_Count12_i_g ;
    wire w_Switch_2;
    wire Game_Inst_o_LED_2_0_i;
    wire w_Switch_4;
    wire Game_Inst_o_LED_4_0_i;
    wire \Game_Inst.N_32 ;
    wire \Game_Inst.N_31 ;
    wire \Game_Inst.r_SM_Main_100_d ;
    wire Game_Inst_o_LED_3_0_i;
    wire \Game_Inst.w_LFSR_Data_9 ;
    wire \Game_Inst.w_LFSR_Data_10 ;
    wire \Game_Inst.w_LFSR_Data_13 ;
    wire \Game_Inst.w_LFSR_Data_14 ;
    wire \Game_Inst.w_LFSR_Data_11 ;
    wire \Game_Inst.w_LFSR_Data_12 ;
    wire \Game_Inst.w_LFSR_Data_15 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_16 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_17 ;
    wire \Game_Inst.LFSR_Inst.r_LFSRZ0Z_18 ;
    wire \Debounce_SW3.r_Count13_10_cascade_ ;
    wire \Debounce_SW3.N_18_2 ;
    wire \Debounce_SW3.N_18_1 ;
    wire \Debounce_SW3.N_18_2_cascade_ ;
    wire \Debounce_SW3.N_20 ;
    wire bfn_11_9_0_;
    wire \Debounce_SW3.r_CountZ0Z_2 ;
    wire \Debounce_SW3.r_Count_1_cry_1 ;
    wire \Debounce_SW3.r_CountZ0Z_3 ;
    wire \Debounce_SW3.r_Count_1_cry_2 ;
    wire \Debounce_SW3.r_CountZ0Z_4 ;
    wire \Debounce_SW3.r_Count_1_cry_3 ;
    wire \Debounce_SW3.r_Count_1_cry_4 ;
    wire \Debounce_SW3.r_CountZ0Z_6 ;
    wire \Debounce_SW3.r_Count_1_cry_5 ;
    wire \Debounce_SW3.r_Count_1_cry_6 ;
    wire \Debounce_SW3.r_CountZ0Z_8 ;
    wire \Debounce_SW3.r_Count_1_cry_7 ;
    wire \Debounce_SW3.r_Count_1_cry_8 ;
    wire \Debounce_SW3.r_CountZ0Z_9 ;
    wire bfn_11_10_0_;
    wire \Debounce_SW3.r_CountZ0Z_10 ;
    wire \Debounce_SW3.r_Count_1_cry_9 ;
    wire \Debounce_SW3.r_CountZ0Z_11 ;
    wire \Debounce_SW3.r_Count_1_cry_10 ;
    wire \Debounce_SW3.r_Count_1_cry_11 ;
    wire \Debounce_SW3.r_Count_1_cry_12 ;
    wire \Debounce_SW3.r_Count_1_cry_13 ;
    wire \Debounce_SW3.r_Count_1_cry_14 ;
    wire \Debounce_SW3.r_Count_1_cry_15 ;
    wire \Debounce_SW3.r_Count_1_cry_16 ;
    wire bfn_11_11_0_;
    wire \Debounce_SW3.r_CountZ0Z_1 ;
    wire \Debounce_SW3.r_CountZ0Z_0 ;
    wire \Debounce_SW3.r_Count12_i_g ;
    wire \Debounce_SW3.N_18 ;
    wire \Debounce_SW3.r_Count12_i ;
    wire \Debounce_SW3.r_CountZ0Z_7 ;
    wire \Debounce_SW3.r_Count13_10 ;
    wire \Debounce_SW3.r_Count13_0_a7_0 ;
    wire \Debounce_SW3.r_Count13_0_a7_4_cascade_ ;
    wire \Debounce_SW3.r_CountZ0Z_5 ;
    wire i_Switch_3_c;
    wire \Debounce_SW3.r_Count13_0_a7_8_cascade_ ;
    wire \Debounce_SW3.r_Count13_0_a7_7 ;
    wire w_Switch_3;
    wire i_Clk_c_g;
    wire \Debounce_SW3.r_CountZ0Z_15 ;
    wire \Debounce_SW3.r_CountZ0Z_13 ;
    wire \Debounce_SW3.r_CountZ0Z_16 ;
    wire \Debounce_SW3.r_CountZ0Z_12 ;
    wire \Debounce_SW3.r_CountZ0Z_17 ;
    wire \Debounce_SW3.un1_r_Count_8lto17_i_2_cascade_ ;
    wire \Debounce_SW3.r_CountZ0Z_14 ;
    wire \Debounce_SW3.un1_r_Count_8lto17_i_3 ;
    wire _gnd_net_;

    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__8737),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__8739),
            .DIN(N__8738),
            .DOUT(N__8737),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__8739),
            .PADOUT(N__8738),
            .PADIN(N__8737),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_4_ibuf_iopad (
            .OE(N__8728),
            .DIN(N__8727),
            .DOUT(N__8726),
            .PACKAGEPIN(i_Switch_4));
    defparam i_Switch_4_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_4_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_4_ibuf_preio (
            .PADOEN(N__8728),
            .PADOUT(N__8727),
            .PADIN(N__8726),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_4_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_1_ibuf_iopad (
            .OE(N__8719),
            .DIN(N__8718),
            .DOUT(N__8717),
            .PACKAGEPIN(i_Switch_1));
    defparam i_Switch_1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_1_ibuf_preio (
            .PADOEN(N__8719),
            .PADOUT(N__8718),
            .PADIN(N__8717),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_3_ibuf_iopad (
            .OE(N__8710),
            .DIN(N__8709),
            .DOUT(N__8708),
            .PACKAGEPIN(i_Switch_3));
    defparam i_Switch_3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_3_ibuf_preio (
            .PADOEN(N__8710),
            .PADOUT(N__8709),
            .PADIN(N__8708),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_2_obuf_iopad (
            .OE(N__8701),
            .DIN(N__8700),
            .DOUT(N__8699),
            .PACKAGEPIN(o_LED_2));
    defparam o_LED_2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_2_obuf_preio (
            .PADOEN(N__8701),
            .PADOUT(N__8700),
            .PADIN(N__8699),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7503),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_E_obuf_iopad (
            .OE(N__8692),
            .DIN(N__8691),
            .DOUT(N__8690),
            .PACKAGEPIN(o_Segment2_E));
    defparam o_Segment2_E_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_E_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_E_obuf_preio (
            .PADOEN(N__8692),
            .PADOUT(N__8691),
            .PADIN(N__8690),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_C_obuf_iopad (
            .OE(N__8683),
            .DIN(N__8682),
            .DOUT(N__8681),
            .PACKAGEPIN(o_Segment2_C));
    defparam o_Segment2_C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_C_obuf_preio (
            .PADOEN(N__8683),
            .PADOUT(N__8682),
            .PADIN(N__8681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4494),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_4_obuf_iopad (
            .OE(N__8674),
            .DIN(N__8673),
            .DOUT(N__8672),
            .PACKAGEPIN(o_LED_4));
    defparam o_LED_4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_4_obuf_preio (
            .PADOEN(N__8674),
            .PADOUT(N__8673),
            .PADIN(N__8672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7452),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_B_obuf_iopad (
            .OE(N__8665),
            .DIN(N__8664),
            .DOUT(N__8663),
            .PACKAGEPIN(o_Segment2_B));
    defparam o_Segment2_B_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_B_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_B_obuf_preio (
            .PADOEN(N__8665),
            .PADOUT(N__8664),
            .PADIN(N__8663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4389),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_3_obuf_iopad (
            .OE(N__8656),
            .DIN(N__8655),
            .DOUT(N__8654),
            .PACKAGEPIN(o_LED_3));
    defparam o_LED_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_3_obuf_preio (
            .PADOEN(N__8656),
            .PADOUT(N__8655),
            .PADIN(N__8654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7836),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_A_obuf_iopad (
            .OE(N__8647),
            .DIN(N__8646),
            .DOUT(N__8645),
            .PACKAGEPIN(o_Segment2_A));
    defparam o_Segment2_A_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_A_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_A_obuf_preio (
            .PADOEN(N__8647),
            .PADOUT(N__8646),
            .PADIN(N__8645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4518),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_G_obuf_iopad (
            .OE(N__8638),
            .DIN(N__8637),
            .DOUT(N__8636),
            .PACKAGEPIN(o_Segment2_G));
    defparam o_Segment2_G_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_G_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_G_obuf_preio (
            .PADOEN(N__8638),
            .PADOUT(N__8637),
            .PADIN(N__8636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4500),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_D_obuf_iopad (
            .OE(N__8629),
            .DIN(N__8628),
            .DOUT(N__8627),
            .PACKAGEPIN(o_Segment2_D));
    defparam o_Segment2_D_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_D_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_D_obuf_preio (
            .PADOEN(N__8629),
            .PADOUT(N__8628),
            .PADIN(N__8627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4506),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_Switch_2_ibuf_iopad (
            .OE(N__8620),
            .DIN(N__8619),
            .DOUT(N__8618),
            .PACKAGEPIN(i_Switch_2));
    defparam i_Switch_2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_Switch_2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Switch_2_ibuf_preio (
            .PADOEN(N__8620),
            .PADOUT(N__8619),
            .PADIN(N__8618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_Switch_2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_Segment2_F_obuf_iopad (
            .OE(N__8611),
            .DIN(N__8610),
            .DOUT(N__8609),
            .PACKAGEPIN(o_Segment2_F));
    defparam o_Segment2_F_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_Segment2_F_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_Segment2_F_obuf_preio (
            .PADOEN(N__8611),
            .PADOUT(N__8610),
            .PADIN(N__8609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4398),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_1_obuf_iopad (
            .OE(N__8602),
            .DIN(N__8601),
            .DOUT(N__8600),
            .PACKAGEPIN(o_LED_1));
    defparam o_LED_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_1_obuf_preio (
            .PADOEN(N__8602),
            .PADOUT(N__8601),
            .PADIN(N__8600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5082),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__1921 (
            .O(N__8583),
            .I(N__8579));
    InMux I__1920 (
            .O(N__8582),
            .I(N__8575));
    InMux I__1919 (
            .O(N__8579),
            .I(N__8572));
    InMux I__1918 (
            .O(N__8578),
            .I(N__8569));
    LocalMux I__1917 (
            .O(N__8575),
            .I(\Debounce_SW3.r_CountZ0Z_7 ));
    LocalMux I__1916 (
            .O(N__8572),
            .I(\Debounce_SW3.r_CountZ0Z_7 ));
    LocalMux I__1915 (
            .O(N__8569),
            .I(\Debounce_SW3.r_CountZ0Z_7 ));
    InMux I__1914 (
            .O(N__8562),
            .I(N__8559));
    LocalMux I__1913 (
            .O(N__8559),
            .I(N__8556));
    Span12Mux_s1_h I__1912 (
            .O(N__8556),
            .I(N__8553));
    Odrv12 I__1911 (
            .O(N__8553),
            .I(\Debounce_SW3.r_Count13_10 ));
    InMux I__1910 (
            .O(N__8550),
            .I(N__8547));
    LocalMux I__1909 (
            .O(N__8547),
            .I(\Debounce_SW3.r_Count13_0_a7_0 ));
    CascadeMux I__1908 (
            .O(N__8544),
            .I(\Debounce_SW3.r_Count13_0_a7_4_cascade_ ));
    InMux I__1907 (
            .O(N__8541),
            .I(N__8536));
    InMux I__1906 (
            .O(N__8540),
            .I(N__8533));
    InMux I__1905 (
            .O(N__8539),
            .I(N__8530));
    LocalMux I__1904 (
            .O(N__8536),
            .I(\Debounce_SW3.r_CountZ0Z_5 ));
    LocalMux I__1903 (
            .O(N__8533),
            .I(\Debounce_SW3.r_CountZ0Z_5 ));
    LocalMux I__1902 (
            .O(N__8530),
            .I(\Debounce_SW3.r_CountZ0Z_5 ));
    CascadeMux I__1901 (
            .O(N__8523),
            .I(N__8519));
    InMux I__1900 (
            .O(N__8522),
            .I(N__8516));
    InMux I__1899 (
            .O(N__8519),
            .I(N__8513));
    LocalMux I__1898 (
            .O(N__8516),
            .I(N__8508));
    LocalMux I__1897 (
            .O(N__8513),
            .I(N__8508));
    Span12Mux_s10_v I__1896 (
            .O(N__8508),
            .I(N__8505));
    Odrv12 I__1895 (
            .O(N__8505),
            .I(i_Switch_3_c));
    CascadeMux I__1894 (
            .O(N__8502),
            .I(\Debounce_SW3.r_Count13_0_a7_8_cascade_ ));
    InMux I__1893 (
            .O(N__8499),
            .I(N__8496));
    LocalMux I__1892 (
            .O(N__8496),
            .I(N__8493));
    Odrv4 I__1891 (
            .O(N__8493),
            .I(\Debounce_SW3.r_Count13_0_a7_7 ));
    InMux I__1890 (
            .O(N__8490),
            .I(N__8486));
    CascadeMux I__1889 (
            .O(N__8489),
            .I(N__8482));
    LocalMux I__1888 (
            .O(N__8486),
            .I(N__8479));
    InMux I__1887 (
            .O(N__8485),
            .I(N__8472));
    InMux I__1886 (
            .O(N__8482),
            .I(N__8472));
    Span4Mux_v I__1885 (
            .O(N__8479),
            .I(N__8469));
    InMux I__1884 (
            .O(N__8478),
            .I(N__8466));
    InMux I__1883 (
            .O(N__8477),
            .I(N__8463));
    LocalMux I__1882 (
            .O(N__8472),
            .I(N__8460));
    Odrv4 I__1881 (
            .O(N__8469),
            .I(w_Switch_3));
    LocalMux I__1880 (
            .O(N__8466),
            .I(w_Switch_3));
    LocalMux I__1879 (
            .O(N__8463),
            .I(w_Switch_3));
    Odrv12 I__1878 (
            .O(N__8460),
            .I(w_Switch_3));
    ClkMux I__1877 (
            .O(N__8451),
            .I(N__8307));
    ClkMux I__1876 (
            .O(N__8450),
            .I(N__8307));
    ClkMux I__1875 (
            .O(N__8449),
            .I(N__8307));
    ClkMux I__1874 (
            .O(N__8448),
            .I(N__8307));
    ClkMux I__1873 (
            .O(N__8447),
            .I(N__8307));
    ClkMux I__1872 (
            .O(N__8446),
            .I(N__8307));
    ClkMux I__1871 (
            .O(N__8445),
            .I(N__8307));
    ClkMux I__1870 (
            .O(N__8444),
            .I(N__8307));
    ClkMux I__1869 (
            .O(N__8443),
            .I(N__8307));
    ClkMux I__1868 (
            .O(N__8442),
            .I(N__8307));
    ClkMux I__1867 (
            .O(N__8441),
            .I(N__8307));
    ClkMux I__1866 (
            .O(N__8440),
            .I(N__8307));
    ClkMux I__1865 (
            .O(N__8439),
            .I(N__8307));
    ClkMux I__1864 (
            .O(N__8438),
            .I(N__8307));
    ClkMux I__1863 (
            .O(N__8437),
            .I(N__8307));
    ClkMux I__1862 (
            .O(N__8436),
            .I(N__8307));
    ClkMux I__1861 (
            .O(N__8435),
            .I(N__8307));
    ClkMux I__1860 (
            .O(N__8434),
            .I(N__8307));
    ClkMux I__1859 (
            .O(N__8433),
            .I(N__8307));
    ClkMux I__1858 (
            .O(N__8432),
            .I(N__8307));
    ClkMux I__1857 (
            .O(N__8431),
            .I(N__8307));
    ClkMux I__1856 (
            .O(N__8430),
            .I(N__8307));
    ClkMux I__1855 (
            .O(N__8429),
            .I(N__8307));
    ClkMux I__1854 (
            .O(N__8428),
            .I(N__8307));
    ClkMux I__1853 (
            .O(N__8427),
            .I(N__8307));
    ClkMux I__1852 (
            .O(N__8426),
            .I(N__8307));
    ClkMux I__1851 (
            .O(N__8425),
            .I(N__8307));
    ClkMux I__1850 (
            .O(N__8424),
            .I(N__8307));
    ClkMux I__1849 (
            .O(N__8423),
            .I(N__8307));
    ClkMux I__1848 (
            .O(N__8422),
            .I(N__8307));
    ClkMux I__1847 (
            .O(N__8421),
            .I(N__8307));
    ClkMux I__1846 (
            .O(N__8420),
            .I(N__8307));
    ClkMux I__1845 (
            .O(N__8419),
            .I(N__8307));
    ClkMux I__1844 (
            .O(N__8418),
            .I(N__8307));
    ClkMux I__1843 (
            .O(N__8417),
            .I(N__8307));
    ClkMux I__1842 (
            .O(N__8416),
            .I(N__8307));
    ClkMux I__1841 (
            .O(N__8415),
            .I(N__8307));
    ClkMux I__1840 (
            .O(N__8414),
            .I(N__8307));
    ClkMux I__1839 (
            .O(N__8413),
            .I(N__8307));
    ClkMux I__1838 (
            .O(N__8412),
            .I(N__8307));
    ClkMux I__1837 (
            .O(N__8411),
            .I(N__8307));
    ClkMux I__1836 (
            .O(N__8410),
            .I(N__8307));
    ClkMux I__1835 (
            .O(N__8409),
            .I(N__8307));
    ClkMux I__1834 (
            .O(N__8408),
            .I(N__8307));
    ClkMux I__1833 (
            .O(N__8407),
            .I(N__8307));
    ClkMux I__1832 (
            .O(N__8406),
            .I(N__8307));
    ClkMux I__1831 (
            .O(N__8405),
            .I(N__8307));
    ClkMux I__1830 (
            .O(N__8404),
            .I(N__8307));
    GlobalMux I__1829 (
            .O(N__8307),
            .I(N__8304));
    gio2CtrlBuf I__1828 (
            .O(N__8304),
            .I(i_Clk_c_g));
    InMux I__1827 (
            .O(N__8301),
            .I(N__8296));
    InMux I__1826 (
            .O(N__8300),
            .I(N__8291));
    InMux I__1825 (
            .O(N__8299),
            .I(N__8291));
    LocalMux I__1824 (
            .O(N__8296),
            .I(\Debounce_SW3.r_CountZ0Z_15 ));
    LocalMux I__1823 (
            .O(N__8291),
            .I(\Debounce_SW3.r_CountZ0Z_15 ));
    InMux I__1822 (
            .O(N__8286),
            .I(N__8282));
    InMux I__1821 (
            .O(N__8285),
            .I(N__8278));
    LocalMux I__1820 (
            .O(N__8282),
            .I(N__8275));
    InMux I__1819 (
            .O(N__8281),
            .I(N__8272));
    LocalMux I__1818 (
            .O(N__8278),
            .I(\Debounce_SW3.r_CountZ0Z_13 ));
    Odrv4 I__1817 (
            .O(N__8275),
            .I(\Debounce_SW3.r_CountZ0Z_13 ));
    LocalMux I__1816 (
            .O(N__8272),
            .I(\Debounce_SW3.r_CountZ0Z_13 ));
    CascadeMux I__1815 (
            .O(N__8265),
            .I(N__8260));
    InMux I__1814 (
            .O(N__8264),
            .I(N__8257));
    InMux I__1813 (
            .O(N__8263),
            .I(N__8252));
    InMux I__1812 (
            .O(N__8260),
            .I(N__8252));
    LocalMux I__1811 (
            .O(N__8257),
            .I(\Debounce_SW3.r_CountZ0Z_16 ));
    LocalMux I__1810 (
            .O(N__8252),
            .I(\Debounce_SW3.r_CountZ0Z_16 ));
    InMux I__1809 (
            .O(N__8247),
            .I(N__8242));
    InMux I__1808 (
            .O(N__8246),
            .I(N__8237));
    InMux I__1807 (
            .O(N__8245),
            .I(N__8237));
    LocalMux I__1806 (
            .O(N__8242),
            .I(\Debounce_SW3.r_CountZ0Z_12 ));
    LocalMux I__1805 (
            .O(N__8237),
            .I(\Debounce_SW3.r_CountZ0Z_12 ));
    InMux I__1804 (
            .O(N__8232),
            .I(N__8227));
    InMux I__1803 (
            .O(N__8231),
            .I(N__8222));
    InMux I__1802 (
            .O(N__8230),
            .I(N__8222));
    LocalMux I__1801 (
            .O(N__8227),
            .I(\Debounce_SW3.r_CountZ0Z_17 ));
    LocalMux I__1800 (
            .O(N__8222),
            .I(\Debounce_SW3.r_CountZ0Z_17 ));
    CascadeMux I__1799 (
            .O(N__8217),
            .I(\Debounce_SW3.un1_r_Count_8lto17_i_2_cascade_ ));
    InMux I__1798 (
            .O(N__8214),
            .I(N__8209));
    InMux I__1797 (
            .O(N__8213),
            .I(N__8204));
    InMux I__1796 (
            .O(N__8212),
            .I(N__8204));
    LocalMux I__1795 (
            .O(N__8209),
            .I(\Debounce_SW3.r_CountZ0Z_14 ));
    LocalMux I__1794 (
            .O(N__8204),
            .I(\Debounce_SW3.r_CountZ0Z_14 ));
    InMux I__1793 (
            .O(N__8199),
            .I(N__8196));
    LocalMux I__1792 (
            .O(N__8196),
            .I(\Debounce_SW3.un1_r_Count_8lto17_i_3 ));
    InMux I__1791 (
            .O(N__8193),
            .I(\Debounce_SW3.r_Count_1_cry_11 ));
    InMux I__1790 (
            .O(N__8190),
            .I(\Debounce_SW3.r_Count_1_cry_12 ));
    InMux I__1789 (
            .O(N__8187),
            .I(\Debounce_SW3.r_Count_1_cry_13 ));
    InMux I__1788 (
            .O(N__8184),
            .I(\Debounce_SW3.r_Count_1_cry_14 ));
    InMux I__1787 (
            .O(N__8181),
            .I(\Debounce_SW3.r_Count_1_cry_15 ));
    InMux I__1786 (
            .O(N__8178),
            .I(bfn_11_11_0_));
    CascadeMux I__1785 (
            .O(N__8175),
            .I(N__8171));
    InMux I__1784 (
            .O(N__8174),
            .I(N__8167));
    InMux I__1783 (
            .O(N__8171),
            .I(N__8164));
    InMux I__1782 (
            .O(N__8170),
            .I(N__8161));
    LocalMux I__1781 (
            .O(N__8167),
            .I(\Debounce_SW3.r_CountZ0Z_1 ));
    LocalMux I__1780 (
            .O(N__8164),
            .I(\Debounce_SW3.r_CountZ0Z_1 ));
    LocalMux I__1779 (
            .O(N__8161),
            .I(\Debounce_SW3.r_CountZ0Z_1 ));
    InMux I__1778 (
            .O(N__8154),
            .I(N__8146));
    InMux I__1777 (
            .O(N__8153),
            .I(N__8146));
    InMux I__1776 (
            .O(N__8152),
            .I(N__8143));
    InMux I__1775 (
            .O(N__8151),
            .I(N__8140));
    LocalMux I__1774 (
            .O(N__8146),
            .I(\Debounce_SW3.r_CountZ0Z_0 ));
    LocalMux I__1773 (
            .O(N__8143),
            .I(\Debounce_SW3.r_CountZ0Z_0 ));
    LocalMux I__1772 (
            .O(N__8140),
            .I(\Debounce_SW3.r_CountZ0Z_0 ));
    SRMux I__1771 (
            .O(N__8133),
            .I(N__8121));
    SRMux I__1770 (
            .O(N__8132),
            .I(N__8121));
    SRMux I__1769 (
            .O(N__8131),
            .I(N__8121));
    SRMux I__1768 (
            .O(N__8130),
            .I(N__8121));
    GlobalMux I__1767 (
            .O(N__8121),
            .I(N__8118));
    gio2CtrlBuf I__1766 (
            .O(N__8118),
            .I(\Debounce_SW3.r_Count12_i_g ));
    InMux I__1765 (
            .O(N__8115),
            .I(N__8112));
    LocalMux I__1764 (
            .O(N__8112),
            .I(\Debounce_SW3.N_18 ));
    IoInMux I__1763 (
            .O(N__8109),
            .I(N__8106));
    LocalMux I__1762 (
            .O(N__8106),
            .I(\Debounce_SW3.r_Count12_i ));
    CascadeMux I__1761 (
            .O(N__8103),
            .I(N__8099));
    InMux I__1760 (
            .O(N__8102),
            .I(N__8096));
    InMux I__1759 (
            .O(N__8099),
            .I(N__8093));
    LocalMux I__1758 (
            .O(N__8096),
            .I(\Debounce_SW3.r_CountZ0Z_3 ));
    LocalMux I__1757 (
            .O(N__8093),
            .I(\Debounce_SW3.r_CountZ0Z_3 ));
    InMux I__1756 (
            .O(N__8088),
            .I(\Debounce_SW3.r_Count_1_cry_2 ));
    InMux I__1755 (
            .O(N__8085),
            .I(N__8080));
    InMux I__1754 (
            .O(N__8084),
            .I(N__8075));
    InMux I__1753 (
            .O(N__8083),
            .I(N__8075));
    LocalMux I__1752 (
            .O(N__8080),
            .I(\Debounce_SW3.r_CountZ0Z_4 ));
    LocalMux I__1751 (
            .O(N__8075),
            .I(\Debounce_SW3.r_CountZ0Z_4 ));
    InMux I__1750 (
            .O(N__8070),
            .I(\Debounce_SW3.r_Count_1_cry_3 ));
    InMux I__1749 (
            .O(N__8067),
            .I(\Debounce_SW3.r_Count_1_cry_4 ));
    InMux I__1748 (
            .O(N__8064),
            .I(N__8059));
    InMux I__1747 (
            .O(N__8063),
            .I(N__8054));
    InMux I__1746 (
            .O(N__8062),
            .I(N__8054));
    LocalMux I__1745 (
            .O(N__8059),
            .I(\Debounce_SW3.r_CountZ0Z_6 ));
    LocalMux I__1744 (
            .O(N__8054),
            .I(\Debounce_SW3.r_CountZ0Z_6 ));
    InMux I__1743 (
            .O(N__8049),
            .I(\Debounce_SW3.r_Count_1_cry_5 ));
    InMux I__1742 (
            .O(N__8046),
            .I(\Debounce_SW3.r_Count_1_cry_6 ));
    InMux I__1741 (
            .O(N__8043),
            .I(N__8039));
    InMux I__1740 (
            .O(N__8042),
            .I(N__8036));
    LocalMux I__1739 (
            .O(N__8039),
            .I(\Debounce_SW3.r_CountZ0Z_8 ));
    LocalMux I__1738 (
            .O(N__8036),
            .I(\Debounce_SW3.r_CountZ0Z_8 ));
    InMux I__1737 (
            .O(N__8031),
            .I(\Debounce_SW3.r_Count_1_cry_7 ));
    InMux I__1736 (
            .O(N__8028),
            .I(N__8024));
    InMux I__1735 (
            .O(N__8027),
            .I(N__8021));
    LocalMux I__1734 (
            .O(N__8024),
            .I(N__8018));
    LocalMux I__1733 (
            .O(N__8021),
            .I(\Debounce_SW3.r_CountZ0Z_9 ));
    Odrv4 I__1732 (
            .O(N__8018),
            .I(\Debounce_SW3.r_CountZ0Z_9 ));
    InMux I__1731 (
            .O(N__8013),
            .I(bfn_11_10_0_));
    InMux I__1730 (
            .O(N__8010),
            .I(N__8006));
    InMux I__1729 (
            .O(N__8009),
            .I(N__8003));
    LocalMux I__1728 (
            .O(N__8006),
            .I(N__8000));
    LocalMux I__1727 (
            .O(N__8003),
            .I(\Debounce_SW3.r_CountZ0Z_10 ));
    Odrv4 I__1726 (
            .O(N__8000),
            .I(\Debounce_SW3.r_CountZ0Z_10 ));
    InMux I__1725 (
            .O(N__7995),
            .I(\Debounce_SW3.r_Count_1_cry_9 ));
    InMux I__1724 (
            .O(N__7992),
            .I(N__7988));
    InMux I__1723 (
            .O(N__7991),
            .I(N__7985));
    LocalMux I__1722 (
            .O(N__7988),
            .I(N__7982));
    LocalMux I__1721 (
            .O(N__7985),
            .I(\Debounce_SW3.r_CountZ0Z_11 ));
    Odrv4 I__1720 (
            .O(N__7982),
            .I(\Debounce_SW3.r_CountZ0Z_11 ));
    InMux I__1719 (
            .O(N__7977),
            .I(\Debounce_SW3.r_Count_1_cry_10 ));
    InMux I__1718 (
            .O(N__7974),
            .I(N__7971));
    LocalMux I__1717 (
            .O(N__7971),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_17 ));
    InMux I__1716 (
            .O(N__7968),
            .I(N__7965));
    LocalMux I__1715 (
            .O(N__7965),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_18 ));
    CascadeMux I__1714 (
            .O(N__7962),
            .I(\Debounce_SW3.r_Count13_10_cascade_ ));
    CascadeMux I__1713 (
            .O(N__7959),
            .I(N__7956));
    InMux I__1712 (
            .O(N__7956),
            .I(N__7953));
    LocalMux I__1711 (
            .O(N__7953),
            .I(\Debounce_SW3.N_18_2 ));
    InMux I__1710 (
            .O(N__7950),
            .I(N__7944));
    InMux I__1709 (
            .O(N__7949),
            .I(N__7944));
    LocalMux I__1708 (
            .O(N__7944),
            .I(\Debounce_SW3.N_18_1 ));
    CascadeMux I__1707 (
            .O(N__7941),
            .I(\Debounce_SW3.N_18_2_cascade_ ));
    InMux I__1706 (
            .O(N__7938),
            .I(N__7935));
    LocalMux I__1705 (
            .O(N__7935),
            .I(\Debounce_SW3.N_20 ));
    InMux I__1704 (
            .O(N__7932),
            .I(N__7928));
    InMux I__1703 (
            .O(N__7931),
            .I(N__7925));
    LocalMux I__1702 (
            .O(N__7928),
            .I(\Debounce_SW3.r_CountZ0Z_2 ));
    LocalMux I__1701 (
            .O(N__7925),
            .I(\Debounce_SW3.r_CountZ0Z_2 ));
    InMux I__1700 (
            .O(N__7920),
            .I(\Debounce_SW3.r_Count_1_cry_1 ));
    InMux I__1699 (
            .O(N__7917),
            .I(N__7908));
    InMux I__1698 (
            .O(N__7916),
            .I(N__7908));
    InMux I__1697 (
            .O(N__7915),
            .I(N__7908));
    LocalMux I__1696 (
            .O(N__7908),
            .I(N__7904));
    InMux I__1695 (
            .O(N__7907),
            .I(N__7901));
    Span4Mux_v I__1694 (
            .O(N__7904),
            .I(N__7897));
    LocalMux I__1693 (
            .O(N__7901),
            .I(N__7894));
    InMux I__1692 (
            .O(N__7900),
            .I(N__7891));
    Odrv4 I__1691 (
            .O(N__7897),
            .I(\Game_Inst.N_32 ));
    Odrv4 I__1690 (
            .O(N__7894),
            .I(\Game_Inst.N_32 ));
    LocalMux I__1689 (
            .O(N__7891),
            .I(\Game_Inst.N_32 ));
    InMux I__1688 (
            .O(N__7884),
            .I(N__7875));
    InMux I__1687 (
            .O(N__7883),
            .I(N__7875));
    InMux I__1686 (
            .O(N__7882),
            .I(N__7875));
    LocalMux I__1685 (
            .O(N__7875),
            .I(N__7871));
    InMux I__1684 (
            .O(N__7874),
            .I(N__7868));
    Span4Mux_v I__1683 (
            .O(N__7871),
            .I(N__7865));
    LocalMux I__1682 (
            .O(N__7868),
            .I(N__7862));
    Odrv4 I__1681 (
            .O(N__7865),
            .I(\Game_Inst.N_31 ));
    Odrv4 I__1680 (
            .O(N__7862),
            .I(\Game_Inst.N_31 ));
    CascadeMux I__1679 (
            .O(N__7857),
            .I(N__7852));
    CascadeMux I__1678 (
            .O(N__7856),
            .I(N__7849));
    InMux I__1677 (
            .O(N__7855),
            .I(N__7842));
    InMux I__1676 (
            .O(N__7852),
            .I(N__7842));
    InMux I__1675 (
            .O(N__7849),
            .I(N__7842));
    LocalMux I__1674 (
            .O(N__7842),
            .I(N__7839));
    Odrv12 I__1673 (
            .O(N__7839),
            .I(\Game_Inst.r_SM_Main_100_d ));
    IoInMux I__1672 (
            .O(N__7836),
            .I(N__7833));
    LocalMux I__1671 (
            .O(N__7833),
            .I(N__7830));
    Odrv4 I__1670 (
            .O(N__7830),
            .I(Game_Inst_o_LED_3_0_i));
    InMux I__1669 (
            .O(N__7827),
            .I(N__7823));
    InMux I__1668 (
            .O(N__7826),
            .I(N__7820));
    LocalMux I__1667 (
            .O(N__7823),
            .I(\Game_Inst.w_LFSR_Data_9 ));
    LocalMux I__1666 (
            .O(N__7820),
            .I(\Game_Inst.w_LFSR_Data_9 ));
    InMux I__1665 (
            .O(N__7815),
            .I(N__7811));
    InMux I__1664 (
            .O(N__7814),
            .I(N__7808));
    LocalMux I__1663 (
            .O(N__7811),
            .I(\Game_Inst.w_LFSR_Data_10 ));
    LocalMux I__1662 (
            .O(N__7808),
            .I(\Game_Inst.w_LFSR_Data_10 ));
    InMux I__1661 (
            .O(N__7803),
            .I(N__7799));
    InMux I__1660 (
            .O(N__7802),
            .I(N__7796));
    LocalMux I__1659 (
            .O(N__7799),
            .I(\Game_Inst.w_LFSR_Data_13 ));
    LocalMux I__1658 (
            .O(N__7796),
            .I(\Game_Inst.w_LFSR_Data_13 ));
    InMux I__1657 (
            .O(N__7791),
            .I(N__7787));
    InMux I__1656 (
            .O(N__7790),
            .I(N__7784));
    LocalMux I__1655 (
            .O(N__7787),
            .I(\Game_Inst.w_LFSR_Data_14 ));
    LocalMux I__1654 (
            .O(N__7784),
            .I(\Game_Inst.w_LFSR_Data_14 ));
    InMux I__1653 (
            .O(N__7779),
            .I(N__7775));
    InMux I__1652 (
            .O(N__7778),
            .I(N__7772));
    LocalMux I__1651 (
            .O(N__7775),
            .I(\Game_Inst.w_LFSR_Data_11 ));
    LocalMux I__1650 (
            .O(N__7772),
            .I(\Game_Inst.w_LFSR_Data_11 ));
    InMux I__1649 (
            .O(N__7767),
            .I(N__7763));
    InMux I__1648 (
            .O(N__7766),
            .I(N__7760));
    LocalMux I__1647 (
            .O(N__7763),
            .I(\Game_Inst.w_LFSR_Data_12 ));
    LocalMux I__1646 (
            .O(N__7760),
            .I(\Game_Inst.w_LFSR_Data_12 ));
    InMux I__1645 (
            .O(N__7755),
            .I(N__7751));
    InMux I__1644 (
            .O(N__7754),
            .I(N__7748));
    LocalMux I__1643 (
            .O(N__7751),
            .I(\Game_Inst.w_LFSR_Data_15 ));
    LocalMux I__1642 (
            .O(N__7748),
            .I(\Game_Inst.w_LFSR_Data_15 ));
    InMux I__1641 (
            .O(N__7743),
            .I(N__7740));
    LocalMux I__1640 (
            .O(N__7740),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_16 ));
    InMux I__1639 (
            .O(N__7737),
            .I(N__7734));
    LocalMux I__1638 (
            .O(N__7734),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_19 ));
    InMux I__1637 (
            .O(N__7731),
            .I(N__7728));
    LocalMux I__1636 (
            .O(N__7728),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_21 ));
    InMux I__1635 (
            .O(N__7725),
            .I(N__7719));
    InMux I__1634 (
            .O(N__7724),
            .I(N__7719));
    LocalMux I__1633 (
            .O(N__7719),
            .I(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_20 ));
    InMux I__1632 (
            .O(N__7716),
            .I(N__7712));
    InMux I__1631 (
            .O(N__7715),
            .I(N__7709));
    LocalMux I__1630 (
            .O(N__7712),
            .I(N__7706));
    LocalMux I__1629 (
            .O(N__7709),
            .I(N__7703));
    Span4Mux_v I__1628 (
            .O(N__7706),
            .I(N__7698));
    Span4Mux_h I__1627 (
            .O(N__7703),
            .I(N__7698));
    Odrv4 I__1626 (
            .O(N__7698),
            .I(\Game_Inst.w_LFSR_Data_0 ));
    InMux I__1625 (
            .O(N__7695),
            .I(N__7690));
    InMux I__1624 (
            .O(N__7694),
            .I(N__7684));
    InMux I__1623 (
            .O(N__7693),
            .I(N__7684));
    LocalMux I__1622 (
            .O(N__7690),
            .I(N__7681));
    InMux I__1621 (
            .O(N__7689),
            .I(N__7678));
    LocalMux I__1620 (
            .O(N__7684),
            .I(\Debounce_SW2.r_CountZ0Z_0 ));
    Odrv4 I__1619 (
            .O(N__7681),
            .I(\Debounce_SW2.r_CountZ0Z_0 ));
    LocalMux I__1618 (
            .O(N__7678),
            .I(\Debounce_SW2.r_CountZ0Z_0 ));
    CascadeMux I__1617 (
            .O(N__7671),
            .I(N__7668));
    InMux I__1616 (
            .O(N__7668),
            .I(N__7664));
    InMux I__1615 (
            .O(N__7667),
            .I(N__7660));
    LocalMux I__1614 (
            .O(N__7664),
            .I(N__7657));
    InMux I__1613 (
            .O(N__7663),
            .I(N__7654));
    LocalMux I__1612 (
            .O(N__7660),
            .I(\Debounce_SW2.r_CountZ0Z_1 ));
    Odrv4 I__1611 (
            .O(N__7657),
            .I(\Debounce_SW2.r_CountZ0Z_1 ));
    LocalMux I__1610 (
            .O(N__7654),
            .I(\Debounce_SW2.r_CountZ0Z_1 ));
    SRMux I__1609 (
            .O(N__7647),
            .I(N__7635));
    SRMux I__1608 (
            .O(N__7646),
            .I(N__7635));
    SRMux I__1607 (
            .O(N__7645),
            .I(N__7635));
    SRMux I__1606 (
            .O(N__7644),
            .I(N__7635));
    GlobalMux I__1605 (
            .O(N__7635),
            .I(N__7632));
    gio2CtrlBuf I__1604 (
            .O(N__7632),
            .I(\Debounce_SW2.r_Count12_i_g ));
    InMux I__1603 (
            .O(N__7629),
            .I(N__7623));
    InMux I__1602 (
            .O(N__7628),
            .I(N__7620));
    InMux I__1601 (
            .O(N__7627),
            .I(N__7617));
    InMux I__1600 (
            .O(N__7626),
            .I(N__7614));
    LocalMux I__1599 (
            .O(N__7623),
            .I(\Debounce_SW4.r_CountZ0Z_0 ));
    LocalMux I__1598 (
            .O(N__7620),
            .I(\Debounce_SW4.r_CountZ0Z_0 ));
    LocalMux I__1597 (
            .O(N__7617),
            .I(\Debounce_SW4.r_CountZ0Z_0 ));
    LocalMux I__1596 (
            .O(N__7614),
            .I(\Debounce_SW4.r_CountZ0Z_0 ));
    SRMux I__1595 (
            .O(N__7605),
            .I(N__7590));
    SRMux I__1594 (
            .O(N__7604),
            .I(N__7590));
    SRMux I__1593 (
            .O(N__7603),
            .I(N__7590));
    SRMux I__1592 (
            .O(N__7602),
            .I(N__7590));
    SRMux I__1591 (
            .O(N__7601),
            .I(N__7590));
    GlobalMux I__1590 (
            .O(N__7590),
            .I(N__7587));
    gio2CtrlBuf I__1589 (
            .O(N__7587),
            .I(\Debounce_SW4.r_Count12_i_g ));
    InMux I__1588 (
            .O(N__7584),
            .I(N__7578));
    InMux I__1587 (
            .O(N__7583),
            .I(N__7574));
    InMux I__1586 (
            .O(N__7582),
            .I(N__7571));
    InMux I__1585 (
            .O(N__7581),
            .I(N__7568));
    LocalMux I__1584 (
            .O(N__7578),
            .I(N__7563));
    InMux I__1583 (
            .O(N__7577),
            .I(N__7560));
    LocalMux I__1582 (
            .O(N__7574),
            .I(N__7557));
    LocalMux I__1581 (
            .O(N__7571),
            .I(N__7552));
    LocalMux I__1580 (
            .O(N__7568),
            .I(N__7549));
    InMux I__1579 (
            .O(N__7567),
            .I(N__7545));
    InMux I__1578 (
            .O(N__7566),
            .I(N__7542));
    Span4Mux_v I__1577 (
            .O(N__7563),
            .I(N__7539));
    LocalMux I__1576 (
            .O(N__7560),
            .I(N__7536));
    Span4Mux_h I__1575 (
            .O(N__7557),
            .I(N__7533));
    InMux I__1574 (
            .O(N__7556),
            .I(N__7528));
    InMux I__1573 (
            .O(N__7555),
            .I(N__7528));
    Span4Mux_h I__1572 (
            .O(N__7552),
            .I(N__7523));
    Span4Mux_h I__1571 (
            .O(N__7549),
            .I(N__7523));
    InMux I__1570 (
            .O(N__7548),
            .I(N__7520));
    LocalMux I__1569 (
            .O(N__7545),
            .I(w_Switch_2));
    LocalMux I__1568 (
            .O(N__7542),
            .I(w_Switch_2));
    Odrv4 I__1567 (
            .O(N__7539),
            .I(w_Switch_2));
    Odrv4 I__1566 (
            .O(N__7536),
            .I(w_Switch_2));
    Odrv4 I__1565 (
            .O(N__7533),
            .I(w_Switch_2));
    LocalMux I__1564 (
            .O(N__7528),
            .I(w_Switch_2));
    Odrv4 I__1563 (
            .O(N__7523),
            .I(w_Switch_2));
    LocalMux I__1562 (
            .O(N__7520),
            .I(w_Switch_2));
    IoInMux I__1561 (
            .O(N__7503),
            .I(N__7500));
    LocalMux I__1560 (
            .O(N__7500),
            .I(N__7497));
    Odrv4 I__1559 (
            .O(N__7497),
            .I(Game_Inst_o_LED_2_0_i));
    CascadeMux I__1558 (
            .O(N__7494),
            .I(N__7491));
    InMux I__1557 (
            .O(N__7491),
            .I(N__7486));
    InMux I__1556 (
            .O(N__7490),
            .I(N__7481));
    InMux I__1555 (
            .O(N__7489),
            .I(N__7481));
    LocalMux I__1554 (
            .O(N__7486),
            .I(N__7478));
    LocalMux I__1553 (
            .O(N__7481),
            .I(N__7473));
    Span4Mux_v I__1552 (
            .O(N__7478),
            .I(N__7470));
    InMux I__1551 (
            .O(N__7477),
            .I(N__7467));
    InMux I__1550 (
            .O(N__7476),
            .I(N__7464));
    Span4Mux_v I__1549 (
            .O(N__7473),
            .I(N__7461));
    Odrv4 I__1548 (
            .O(N__7470),
            .I(w_Switch_4));
    LocalMux I__1547 (
            .O(N__7467),
            .I(w_Switch_4));
    LocalMux I__1546 (
            .O(N__7464),
            .I(w_Switch_4));
    Odrv4 I__1545 (
            .O(N__7461),
            .I(w_Switch_4));
    IoInMux I__1544 (
            .O(N__7452),
            .I(N__7449));
    LocalMux I__1543 (
            .O(N__7449),
            .I(N__7446));
    Span4Mux_s3_h I__1542 (
            .O(N__7446),
            .I(N__7443));
    Odrv4 I__1541 (
            .O(N__7443),
            .I(Game_Inst_o_LED_4_0_i));
    InMux I__1540 (
            .O(N__7440),
            .I(N__7437));
    LocalMux I__1539 (
            .O(N__7437),
            .I(\Game_Inst.r_Pattern_5_Z0Z_0 ));
    InMux I__1538 (
            .O(N__7434),
            .I(N__7431));
    LocalMux I__1537 (
            .O(N__7431),
            .I(N__7428));
    Odrv4 I__1536 (
            .O(N__7428),
            .I(\Game_Inst.r_Pattern_5_Z0Z_1 ));
    InMux I__1535 (
            .O(N__7425),
            .I(N__7422));
    LocalMux I__1534 (
            .O(N__7422),
            .I(\Game_Inst.r_Pattern_6_Z0Z_0 ));
    InMux I__1533 (
            .O(N__7419),
            .I(N__7416));
    LocalMux I__1532 (
            .O(N__7416),
            .I(\Game_Inst.r_Pattern_6_Z0Z_1 ));
    InMux I__1531 (
            .O(N__7413),
            .I(N__7410));
    LocalMux I__1530 (
            .O(N__7410),
            .I(\Game_Inst.r_Pattern_7_Z0Z_0 ));
    InMux I__1529 (
            .O(N__7407),
            .I(N__7404));
    LocalMux I__1528 (
            .O(N__7404),
            .I(\Game_Inst.r_Pattern_7_Z0Z_1 ));
    CEMux I__1527 (
            .O(N__7401),
            .I(N__7397));
    CEMux I__1526 (
            .O(N__7400),
            .I(N__7394));
    LocalMux I__1525 (
            .O(N__7397),
            .I(N__7390));
    LocalMux I__1524 (
            .O(N__7394),
            .I(N__7387));
    CEMux I__1523 (
            .O(N__7393),
            .I(N__7384));
    Span4Mux_h I__1522 (
            .O(N__7390),
            .I(N__7381));
    Span4Mux_h I__1521 (
            .O(N__7387),
            .I(N__7378));
    LocalMux I__1520 (
            .O(N__7384),
            .I(N__7375));
    Span4Mux_h I__1519 (
            .O(N__7381),
            .I(N__7372));
    Span4Mux_h I__1518 (
            .O(N__7378),
            .I(N__7369));
    Span4Mux_h I__1517 (
            .O(N__7375),
            .I(N__7366));
    Odrv4 I__1516 (
            .O(N__7372),
            .I(\Game_Inst.r_SM_Main_98_d ));
    Odrv4 I__1515 (
            .O(N__7369),
            .I(\Game_Inst.r_SM_Main_98_d ));
    Odrv4 I__1514 (
            .O(N__7366),
            .I(\Game_Inst.r_SM_Main_98_d ));
    InMux I__1513 (
            .O(N__7359),
            .I(N__7355));
    InMux I__1512 (
            .O(N__7358),
            .I(N__7352));
    LocalMux I__1511 (
            .O(N__7355),
            .I(N__7349));
    LocalMux I__1510 (
            .O(N__7352),
            .I(N__7345));
    Span12Mux_s9_v I__1509 (
            .O(N__7349),
            .I(N__7342));
    InMux I__1508 (
            .O(N__7348),
            .I(N__7339));
    Odrv4 I__1507 (
            .O(N__7345),
            .I(\Game_Inst.r_Button_ID_2_sm0_0 ));
    Odrv12 I__1506 (
            .O(N__7342),
            .I(\Game_Inst.r_Button_ID_2_sm0_0 ));
    LocalMux I__1505 (
            .O(N__7339),
            .I(\Game_Inst.r_Button_ID_2_sm0_0 ));
    InMux I__1504 (
            .O(N__7332),
            .I(N__7328));
    InMux I__1503 (
            .O(N__7331),
            .I(N__7325));
    LocalMux I__1502 (
            .O(N__7328),
            .I(\Game_Inst.r_SwitchZ0Z_2 ));
    LocalMux I__1501 (
            .O(N__7325),
            .I(\Game_Inst.r_SwitchZ0Z_2 ));
    InMux I__1500 (
            .O(N__7320),
            .I(N__7317));
    LocalMux I__1499 (
            .O(N__7317),
            .I(\Game_Inst.r_SwitchZ0Z_3 ));
    InMux I__1498 (
            .O(N__7314),
            .I(\Debounce_SW4.r_Count_1_cry_14 ));
    InMux I__1497 (
            .O(N__7311),
            .I(N__7306));
    InMux I__1496 (
            .O(N__7310),
            .I(N__7301));
    InMux I__1495 (
            .O(N__7309),
            .I(N__7301));
    LocalMux I__1494 (
            .O(N__7306),
            .I(\Debounce_SW4.r_CountZ0Z_16 ));
    LocalMux I__1493 (
            .O(N__7301),
            .I(\Debounce_SW4.r_CountZ0Z_16 ));
    InMux I__1492 (
            .O(N__7296),
            .I(\Debounce_SW4.r_Count_1_cry_15 ));
    InMux I__1491 (
            .O(N__7293),
            .I(bfn_8_7_0_));
    CascadeMux I__1490 (
            .O(N__7290),
            .I(N__7285));
    CascadeMux I__1489 (
            .O(N__7289),
            .I(N__7282));
    InMux I__1488 (
            .O(N__7288),
            .I(N__7279));
    InMux I__1487 (
            .O(N__7285),
            .I(N__7274));
    InMux I__1486 (
            .O(N__7282),
            .I(N__7274));
    LocalMux I__1485 (
            .O(N__7279),
            .I(\Debounce_SW4.r_CountZ0Z_17 ));
    LocalMux I__1484 (
            .O(N__7274),
            .I(\Debounce_SW4.r_CountZ0Z_17 ));
    InMux I__1483 (
            .O(N__7269),
            .I(N__7265));
    InMux I__1482 (
            .O(N__7268),
            .I(N__7262));
    LocalMux I__1481 (
            .O(N__7265),
            .I(\Game_Inst.w_LFSR_Data_7 ));
    LocalMux I__1480 (
            .O(N__7262),
            .I(\Game_Inst.w_LFSR_Data_7 ));
    InMux I__1479 (
            .O(N__7257),
            .I(N__7253));
    InMux I__1478 (
            .O(N__7256),
            .I(N__7250));
    LocalMux I__1477 (
            .O(N__7253),
            .I(N__7247));
    LocalMux I__1476 (
            .O(N__7250),
            .I(\Game_Inst.w_LFSR_Data_5 ));
    Odrv4 I__1475 (
            .O(N__7247),
            .I(\Game_Inst.w_LFSR_Data_5 ));
    InMux I__1474 (
            .O(N__7242),
            .I(N__7238));
    InMux I__1473 (
            .O(N__7241),
            .I(N__7235));
    LocalMux I__1472 (
            .O(N__7238),
            .I(\Game_Inst.w_LFSR_Data_6 ));
    LocalMux I__1471 (
            .O(N__7235),
            .I(\Game_Inst.w_LFSR_Data_6 ));
    InMux I__1470 (
            .O(N__7230),
            .I(N__7226));
    InMux I__1469 (
            .O(N__7229),
            .I(N__7223));
    LocalMux I__1468 (
            .O(N__7226),
            .I(\Game_Inst.w_LFSR_Data_8 ));
    LocalMux I__1467 (
            .O(N__7223),
            .I(\Game_Inst.w_LFSR_Data_8 ));
    InMux I__1466 (
            .O(N__7218),
            .I(N__7215));
    LocalMux I__1465 (
            .O(N__7215),
            .I(\Game_Inst.r_Pattern_4_Z0Z_0 ));
    InMux I__1464 (
            .O(N__7212),
            .I(N__7209));
    LocalMux I__1463 (
            .O(N__7209),
            .I(N__7206));
    Odrv4 I__1462 (
            .O(N__7206),
            .I(\Game_Inst.r_Pattern_4_Z0Z_1 ));
    InMux I__1461 (
            .O(N__7203),
            .I(N__7198));
    InMux I__1460 (
            .O(N__7202),
            .I(N__7195));
    InMux I__1459 (
            .O(N__7201),
            .I(N__7192));
    LocalMux I__1458 (
            .O(N__7198),
            .I(\Debounce_SW4.r_CountZ0Z_7 ));
    LocalMux I__1457 (
            .O(N__7195),
            .I(\Debounce_SW4.r_CountZ0Z_7 ));
    LocalMux I__1456 (
            .O(N__7192),
            .I(\Debounce_SW4.r_CountZ0Z_7 ));
    InMux I__1455 (
            .O(N__7185),
            .I(\Debounce_SW4.r_Count_1_cry_6 ));
    InMux I__1454 (
            .O(N__7182),
            .I(N__7177));
    InMux I__1453 (
            .O(N__7181),
            .I(N__7172));
    InMux I__1452 (
            .O(N__7180),
            .I(N__7172));
    LocalMux I__1451 (
            .O(N__7177),
            .I(\Debounce_SW4.r_CountZ0Z_8 ));
    LocalMux I__1450 (
            .O(N__7172),
            .I(\Debounce_SW4.r_CountZ0Z_8 ));
    InMux I__1449 (
            .O(N__7167),
            .I(\Debounce_SW4.r_Count_1_cry_7 ));
    InMux I__1448 (
            .O(N__7164),
            .I(N__7159));
    InMux I__1447 (
            .O(N__7163),
            .I(N__7156));
    InMux I__1446 (
            .O(N__7162),
            .I(N__7153));
    LocalMux I__1445 (
            .O(N__7159),
            .I(\Debounce_SW4.r_CountZ0Z_9 ));
    LocalMux I__1444 (
            .O(N__7156),
            .I(\Debounce_SW4.r_CountZ0Z_9 ));
    LocalMux I__1443 (
            .O(N__7153),
            .I(\Debounce_SW4.r_CountZ0Z_9 ));
    InMux I__1442 (
            .O(N__7146),
            .I(bfn_8_6_0_));
    InMux I__1441 (
            .O(N__7143),
            .I(N__7138));
    InMux I__1440 (
            .O(N__7142),
            .I(N__7133));
    InMux I__1439 (
            .O(N__7141),
            .I(N__7133));
    LocalMux I__1438 (
            .O(N__7138),
            .I(\Debounce_SW4.r_CountZ0Z_10 ));
    LocalMux I__1437 (
            .O(N__7133),
            .I(\Debounce_SW4.r_CountZ0Z_10 ));
    InMux I__1436 (
            .O(N__7128),
            .I(\Debounce_SW4.r_Count_1_cry_9 ));
    CascadeMux I__1435 (
            .O(N__7125),
            .I(N__7120));
    InMux I__1434 (
            .O(N__7124),
            .I(N__7117));
    InMux I__1433 (
            .O(N__7123),
            .I(N__7114));
    InMux I__1432 (
            .O(N__7120),
            .I(N__7111));
    LocalMux I__1431 (
            .O(N__7117),
            .I(\Debounce_SW4.r_CountZ0Z_11 ));
    LocalMux I__1430 (
            .O(N__7114),
            .I(\Debounce_SW4.r_CountZ0Z_11 ));
    LocalMux I__1429 (
            .O(N__7111),
            .I(\Debounce_SW4.r_CountZ0Z_11 ));
    InMux I__1428 (
            .O(N__7104),
            .I(\Debounce_SW4.r_Count_1_cry_10 ));
    InMux I__1427 (
            .O(N__7101),
            .I(N__7096));
    InMux I__1426 (
            .O(N__7100),
            .I(N__7093));
    InMux I__1425 (
            .O(N__7099),
            .I(N__7090));
    LocalMux I__1424 (
            .O(N__7096),
            .I(\Debounce_SW4.r_CountZ0Z_12 ));
    LocalMux I__1423 (
            .O(N__7093),
            .I(\Debounce_SW4.r_CountZ0Z_12 ));
    LocalMux I__1422 (
            .O(N__7090),
            .I(\Debounce_SW4.r_CountZ0Z_12 ));
    InMux I__1421 (
            .O(N__7083),
            .I(\Debounce_SW4.r_Count_1_cry_11 ));
    CascadeMux I__1420 (
            .O(N__7080),
            .I(N__7075));
    InMux I__1419 (
            .O(N__7079),
            .I(N__7072));
    InMux I__1418 (
            .O(N__7078),
            .I(N__7069));
    InMux I__1417 (
            .O(N__7075),
            .I(N__7066));
    LocalMux I__1416 (
            .O(N__7072),
            .I(N__7063));
    LocalMux I__1415 (
            .O(N__7069),
            .I(\Debounce_SW4.r_CountZ0Z_13 ));
    LocalMux I__1414 (
            .O(N__7066),
            .I(\Debounce_SW4.r_CountZ0Z_13 ));
    Odrv4 I__1413 (
            .O(N__7063),
            .I(\Debounce_SW4.r_CountZ0Z_13 ));
    InMux I__1412 (
            .O(N__7056),
            .I(\Debounce_SW4.r_Count_1_cry_12 ));
    InMux I__1411 (
            .O(N__7053),
            .I(N__7048));
    InMux I__1410 (
            .O(N__7052),
            .I(N__7043));
    InMux I__1409 (
            .O(N__7051),
            .I(N__7043));
    LocalMux I__1408 (
            .O(N__7048),
            .I(\Debounce_SW4.r_CountZ0Z_14 ));
    LocalMux I__1407 (
            .O(N__7043),
            .I(\Debounce_SW4.r_CountZ0Z_14 ));
    InMux I__1406 (
            .O(N__7038),
            .I(\Debounce_SW4.r_Count_1_cry_13 ));
    InMux I__1405 (
            .O(N__7035),
            .I(N__7030));
    InMux I__1404 (
            .O(N__7034),
            .I(N__7025));
    InMux I__1403 (
            .O(N__7033),
            .I(N__7025));
    LocalMux I__1402 (
            .O(N__7030),
            .I(\Debounce_SW4.r_CountZ0Z_15 ));
    LocalMux I__1401 (
            .O(N__7025),
            .I(\Debounce_SW4.r_CountZ0Z_15 ));
    InMux I__1400 (
            .O(N__7020),
            .I(N__7015));
    InMux I__1399 (
            .O(N__7019),
            .I(N__7010));
    InMux I__1398 (
            .O(N__7018),
            .I(N__7010));
    LocalMux I__1397 (
            .O(N__7015),
            .I(N__7005));
    LocalMux I__1396 (
            .O(N__7010),
            .I(N__7005));
    Odrv4 I__1395 (
            .O(N__7005),
            .I(\Debounce_SW2.r_CountZ0Z_12 ));
    InMux I__1394 (
            .O(N__7002),
            .I(N__6999));
    LocalMux I__1393 (
            .O(N__6999),
            .I(\Debounce_SW2.r_Count13_0_a7_4 ));
    InMux I__1392 (
            .O(N__6996),
            .I(N__6990));
    InMux I__1391 (
            .O(N__6995),
            .I(N__6990));
    LocalMux I__1390 (
            .O(N__6990),
            .I(\Debounce_SW4.r_Count13_10 ));
    CascadeMux I__1389 (
            .O(N__6987),
            .I(N__6984));
    InMux I__1388 (
            .O(N__6984),
            .I(N__6980));
    InMux I__1387 (
            .O(N__6983),
            .I(N__6976));
    LocalMux I__1386 (
            .O(N__6980),
            .I(N__6973));
    InMux I__1385 (
            .O(N__6979),
            .I(N__6970));
    LocalMux I__1384 (
            .O(N__6976),
            .I(\Debounce_SW4.r_CountZ0Z_1 ));
    Odrv4 I__1383 (
            .O(N__6973),
            .I(\Debounce_SW4.r_CountZ0Z_1 ));
    LocalMux I__1382 (
            .O(N__6970),
            .I(\Debounce_SW4.r_CountZ0Z_1 ));
    InMux I__1381 (
            .O(N__6963),
            .I(N__6959));
    InMux I__1380 (
            .O(N__6962),
            .I(N__6956));
    LocalMux I__1379 (
            .O(N__6959),
            .I(\Debounce_SW4.r_CountZ0Z_2 ));
    LocalMux I__1378 (
            .O(N__6956),
            .I(\Debounce_SW4.r_CountZ0Z_2 ));
    InMux I__1377 (
            .O(N__6951),
            .I(\Debounce_SW4.r_Count_1_cry_1 ));
    CascadeMux I__1376 (
            .O(N__6948),
            .I(N__6944));
    InMux I__1375 (
            .O(N__6947),
            .I(N__6941));
    InMux I__1374 (
            .O(N__6944),
            .I(N__6938));
    LocalMux I__1373 (
            .O(N__6941),
            .I(\Debounce_SW4.r_CountZ0Z_3 ));
    LocalMux I__1372 (
            .O(N__6938),
            .I(\Debounce_SW4.r_CountZ0Z_3 ));
    InMux I__1371 (
            .O(N__6933),
            .I(\Debounce_SW4.r_Count_1_cry_2 ));
    InMux I__1370 (
            .O(N__6930),
            .I(N__6926));
    InMux I__1369 (
            .O(N__6929),
            .I(N__6923));
    LocalMux I__1368 (
            .O(N__6926),
            .I(\Debounce_SW4.r_CountZ0Z_4 ));
    LocalMux I__1367 (
            .O(N__6923),
            .I(\Debounce_SW4.r_CountZ0Z_4 ));
    InMux I__1366 (
            .O(N__6918),
            .I(\Debounce_SW4.r_Count_1_cry_3 ));
    InMux I__1365 (
            .O(N__6915),
            .I(N__6911));
    InMux I__1364 (
            .O(N__6914),
            .I(N__6908));
    LocalMux I__1363 (
            .O(N__6911),
            .I(\Debounce_SW4.r_CountZ0Z_5 ));
    LocalMux I__1362 (
            .O(N__6908),
            .I(\Debounce_SW4.r_CountZ0Z_5 ));
    InMux I__1361 (
            .O(N__6903),
            .I(\Debounce_SW4.r_Count_1_cry_4 ));
    CascadeMux I__1360 (
            .O(N__6900),
            .I(N__6896));
    InMux I__1359 (
            .O(N__6899),
            .I(N__6892));
    InMux I__1358 (
            .O(N__6896),
            .I(N__6887));
    InMux I__1357 (
            .O(N__6895),
            .I(N__6887));
    LocalMux I__1356 (
            .O(N__6892),
            .I(\Debounce_SW4.r_CountZ0Z_6 ));
    LocalMux I__1355 (
            .O(N__6887),
            .I(\Debounce_SW4.r_CountZ0Z_6 ));
    InMux I__1354 (
            .O(N__6882),
            .I(\Debounce_SW4.r_Count_1_cry_5 ));
    InMux I__1353 (
            .O(N__6879),
            .I(N__6875));
    InMux I__1352 (
            .O(N__6878),
            .I(N__6872));
    LocalMux I__1351 (
            .O(N__6875),
            .I(\Debounce_SW2.r_CountZ0Z_8 ));
    LocalMux I__1350 (
            .O(N__6872),
            .I(\Debounce_SW2.r_CountZ0Z_8 ));
    CascadeMux I__1349 (
            .O(N__6867),
            .I(N__6864));
    InMux I__1348 (
            .O(N__6864),
            .I(N__6861));
    LocalMux I__1347 (
            .O(N__6861),
            .I(\Debounce_SW2.r_Count13_10 ));
    InMux I__1346 (
            .O(N__6858),
            .I(N__6853));
    InMux I__1345 (
            .O(N__6857),
            .I(N__6848));
    InMux I__1344 (
            .O(N__6856),
            .I(N__6848));
    LocalMux I__1343 (
            .O(N__6853),
            .I(\Debounce_SW2.r_CountZ0Z_5 ));
    LocalMux I__1342 (
            .O(N__6848),
            .I(\Debounce_SW2.r_CountZ0Z_5 ));
    InMux I__1341 (
            .O(N__6843),
            .I(N__6840));
    LocalMux I__1340 (
            .O(N__6840),
            .I(N__6837));
    Odrv4 I__1339 (
            .O(N__6837),
            .I(\Debounce_SW2.r_Count13_0_a7_8 ));
    InMux I__1338 (
            .O(N__6834),
            .I(N__6831));
    LocalMux I__1337 (
            .O(N__6831),
            .I(\Debounce_SW2.r_Count13_0_a7_0 ));
    InMux I__1336 (
            .O(N__6828),
            .I(N__6824));
    InMux I__1335 (
            .O(N__6827),
            .I(N__6821));
    LocalMux I__1334 (
            .O(N__6824),
            .I(\Debounce_SW2.r_CountZ0Z_9 ));
    LocalMux I__1333 (
            .O(N__6821),
            .I(\Debounce_SW2.r_CountZ0Z_9 ));
    InMux I__1332 (
            .O(N__6816),
            .I(N__6812));
    InMux I__1331 (
            .O(N__6815),
            .I(N__6809));
    LocalMux I__1330 (
            .O(N__6812),
            .I(\Debounce_SW2.r_CountZ0Z_10 ));
    LocalMux I__1329 (
            .O(N__6809),
            .I(\Debounce_SW2.r_CountZ0Z_10 ));
    CascadeMux I__1328 (
            .O(N__6804),
            .I(N__6801));
    InMux I__1327 (
            .O(N__6801),
            .I(N__6798));
    LocalMux I__1326 (
            .O(N__6798),
            .I(N__6795));
    Odrv4 I__1325 (
            .O(N__6795),
            .I(\Debounce_SW2.N_23_2 ));
    InMux I__1324 (
            .O(N__6792),
            .I(N__6788));
    InMux I__1323 (
            .O(N__6791),
            .I(N__6785));
    LocalMux I__1322 (
            .O(N__6788),
            .I(\Debounce_SW2.N_23_1 ));
    LocalMux I__1321 (
            .O(N__6785),
            .I(\Debounce_SW2.N_23_1 ));
    CascadeMux I__1320 (
            .O(N__6780),
            .I(\Debounce_SW2.N_23_2_cascade_ ));
    InMux I__1319 (
            .O(N__6777),
            .I(N__6774));
    LocalMux I__1318 (
            .O(N__6774),
            .I(\Debounce_SW2.N_25 ));
    InMux I__1317 (
            .O(N__6771),
            .I(N__6767));
    CascadeMux I__1316 (
            .O(N__6770),
            .I(N__6764));
    LocalMux I__1315 (
            .O(N__6767),
            .I(N__6761));
    InMux I__1314 (
            .O(N__6764),
            .I(N__6758));
    Span4Mux_v I__1313 (
            .O(N__6761),
            .I(N__6753));
    LocalMux I__1312 (
            .O(N__6758),
            .I(N__6753));
    Span4Mux_v I__1311 (
            .O(N__6753),
            .I(N__6750));
    Span4Mux_h I__1310 (
            .O(N__6750),
            .I(N__6747));
    Span4Mux_v I__1309 (
            .O(N__6747),
            .I(N__6744));
    Odrv4 I__1308 (
            .O(N__6744),
            .I(i_Switch_2_c));
    CascadeMux I__1307 (
            .O(N__6741),
            .I(\Debounce_SW2.N_23_cascade_ ));
    IoInMux I__1306 (
            .O(N__6738),
            .I(N__6735));
    LocalMux I__1305 (
            .O(N__6735),
            .I(N__6732));
    Span4Mux_s2_v I__1304 (
            .O(N__6732),
            .I(N__6729));
    Odrv4 I__1303 (
            .O(N__6729),
            .I(\Debounce_SW2.r_Count12_i ));
    InMux I__1302 (
            .O(N__6726),
            .I(N__6721));
    InMux I__1301 (
            .O(N__6725),
            .I(N__6716));
    InMux I__1300 (
            .O(N__6724),
            .I(N__6716));
    LocalMux I__1299 (
            .O(N__6721),
            .I(\Debounce_SW2.r_CountZ0Z_15 ));
    LocalMux I__1298 (
            .O(N__6716),
            .I(\Debounce_SW2.r_CountZ0Z_15 ));
    InMux I__1297 (
            .O(N__6711),
            .I(N__6706));
    InMux I__1296 (
            .O(N__6710),
            .I(N__6701));
    InMux I__1295 (
            .O(N__6709),
            .I(N__6701));
    LocalMux I__1294 (
            .O(N__6706),
            .I(\Debounce_SW2.r_CountZ0Z_13 ));
    LocalMux I__1293 (
            .O(N__6701),
            .I(\Debounce_SW2.r_CountZ0Z_13 ));
    InMux I__1292 (
            .O(N__6696),
            .I(N__6691));
    InMux I__1291 (
            .O(N__6695),
            .I(N__6686));
    InMux I__1290 (
            .O(N__6694),
            .I(N__6686));
    LocalMux I__1289 (
            .O(N__6691),
            .I(\Debounce_SW2.r_CountZ0Z_14 ));
    LocalMux I__1288 (
            .O(N__6686),
            .I(\Debounce_SW2.r_CountZ0Z_14 ));
    CascadeMux I__1287 (
            .O(N__6681),
            .I(\Debounce_SW2.un1_r_Count_8lto17_i_2_cascade_ ));
    InMux I__1286 (
            .O(N__6678),
            .I(N__6675));
    LocalMux I__1285 (
            .O(N__6675),
            .I(\Debounce_SW2.un1_r_Count_8lto17_i_3 ));
    CascadeMux I__1284 (
            .O(N__6672),
            .I(N__6667));
    InMux I__1283 (
            .O(N__6671),
            .I(N__6664));
    InMux I__1282 (
            .O(N__6670),
            .I(N__6659));
    InMux I__1281 (
            .O(N__6667),
            .I(N__6659));
    LocalMux I__1280 (
            .O(N__6664),
            .I(\Debounce_SW2.r_CountZ0Z_16 ));
    LocalMux I__1279 (
            .O(N__6659),
            .I(\Debounce_SW2.r_CountZ0Z_16 ));
    InMux I__1278 (
            .O(N__6654),
            .I(N__6649));
    InMux I__1277 (
            .O(N__6653),
            .I(N__6646));
    InMux I__1276 (
            .O(N__6652),
            .I(N__6643));
    LocalMux I__1275 (
            .O(N__6649),
            .I(\Debounce_SW2.r_CountZ0Z_17 ));
    LocalMux I__1274 (
            .O(N__6646),
            .I(\Debounce_SW2.r_CountZ0Z_17 ));
    LocalMux I__1273 (
            .O(N__6643),
            .I(\Debounce_SW2.r_CountZ0Z_17 ));
    CascadeMux I__1272 (
            .O(N__6636),
            .I(N__6632));
    InMux I__1271 (
            .O(N__6635),
            .I(N__6628));
    InMux I__1270 (
            .O(N__6632),
            .I(N__6623));
    InMux I__1269 (
            .O(N__6631),
            .I(N__6623));
    LocalMux I__1268 (
            .O(N__6628),
            .I(\Debounce_SW2.r_CountZ0Z_7 ));
    LocalMux I__1267 (
            .O(N__6623),
            .I(\Debounce_SW2.r_CountZ0Z_7 ));
    CascadeMux I__1266 (
            .O(N__6618),
            .I(N__6615));
    InMux I__1265 (
            .O(N__6615),
            .I(N__6612));
    LocalMux I__1264 (
            .O(N__6612),
            .I(\Game_Inst.r_Pattern_6__RNINHCKZ0Z_0 ));
    InMux I__1263 (
            .O(N__6609),
            .I(N__6606));
    LocalMux I__1262 (
            .O(N__6606),
            .I(N__6602));
    InMux I__1261 (
            .O(N__6605),
            .I(N__6599));
    Odrv4 I__1260 (
            .O(N__6602),
            .I(\Game_Inst.w_LFSR_Data_1 ));
    LocalMux I__1259 (
            .O(N__6599),
            .I(\Game_Inst.w_LFSR_Data_1 ));
    InMux I__1258 (
            .O(N__6594),
            .I(N__6590));
    InMux I__1257 (
            .O(N__6593),
            .I(N__6587));
    LocalMux I__1256 (
            .O(N__6590),
            .I(\Game_Inst.w_LFSR_Data_2 ));
    LocalMux I__1255 (
            .O(N__6587),
            .I(\Game_Inst.w_LFSR_Data_2 ));
    CascadeMux I__1254 (
            .O(N__6582),
            .I(N__6579));
    InMux I__1253 (
            .O(N__6579),
            .I(N__6575));
    InMux I__1252 (
            .O(N__6578),
            .I(N__6572));
    LocalMux I__1251 (
            .O(N__6575),
            .I(N__6557));
    LocalMux I__1250 (
            .O(N__6572),
            .I(N__6557));
    InMux I__1249 (
            .O(N__6571),
            .I(N__6554));
    InMux I__1248 (
            .O(N__6570),
            .I(N__6549));
    InMux I__1247 (
            .O(N__6569),
            .I(N__6549));
    InMux I__1246 (
            .O(N__6568),
            .I(N__6542));
    InMux I__1245 (
            .O(N__6567),
            .I(N__6542));
    InMux I__1244 (
            .O(N__6566),
            .I(N__6542));
    InMux I__1243 (
            .O(N__6565),
            .I(N__6537));
    InMux I__1242 (
            .O(N__6564),
            .I(N__6537));
    InMux I__1241 (
            .O(N__6563),
            .I(N__6532));
    InMux I__1240 (
            .O(N__6562),
            .I(N__6532));
    Odrv4 I__1239 (
            .O(N__6557),
            .I(\Game_Inst.r_IndexZ0Z_0 ));
    LocalMux I__1238 (
            .O(N__6554),
            .I(\Game_Inst.r_IndexZ0Z_0 ));
    LocalMux I__1237 (
            .O(N__6549),
            .I(\Game_Inst.r_IndexZ0Z_0 ));
    LocalMux I__1236 (
            .O(N__6542),
            .I(\Game_Inst.r_IndexZ0Z_0 ));
    LocalMux I__1235 (
            .O(N__6537),
            .I(\Game_Inst.r_IndexZ0Z_0 ));
    LocalMux I__1234 (
            .O(N__6532),
            .I(\Game_Inst.r_IndexZ0Z_0 ));
    InMux I__1233 (
            .O(N__6519),
            .I(N__6516));
    LocalMux I__1232 (
            .O(N__6516),
            .I(\Game_Inst.r_Pattern_5__RNIJ1KJZ0Z_0 ));
    InMux I__1231 (
            .O(N__6513),
            .I(N__6510));
    LocalMux I__1230 (
            .O(N__6510),
            .I(N__6506));
    CascadeMux I__1229 (
            .O(N__6509),
            .I(N__6503));
    Span4Mux_v I__1228 (
            .O(N__6506),
            .I(N__6500));
    InMux I__1227 (
            .O(N__6503),
            .I(N__6497));
    Odrv4 I__1226 (
            .O(N__6500),
            .I(\Game_Inst.un1_i_Switch_4_1 ));
    LocalMux I__1225 (
            .O(N__6497),
            .I(\Game_Inst.un1_i_Switch_4_1 ));
    InMux I__1224 (
            .O(N__6492),
            .I(N__6486));
    InMux I__1223 (
            .O(N__6491),
            .I(N__6486));
    LocalMux I__1222 (
            .O(N__6486),
            .I(\Game_Inst.r_Button_ID_2_0 ));
    InMux I__1221 (
            .O(N__6483),
            .I(N__6480));
    LocalMux I__1220 (
            .O(N__6480),
            .I(\Debounce_SW2.r_Count13_0_a7_7 ));
    InMux I__1219 (
            .O(N__6477),
            .I(N__6473));
    InMux I__1218 (
            .O(N__6476),
            .I(N__6470));
    LocalMux I__1217 (
            .O(N__6473),
            .I(\Debounce_SW2.r_CountZ0Z_2 ));
    LocalMux I__1216 (
            .O(N__6470),
            .I(\Debounce_SW2.r_CountZ0Z_2 ));
    CascadeMux I__1215 (
            .O(N__6465),
            .I(N__6461));
    InMux I__1214 (
            .O(N__6464),
            .I(N__6458));
    InMux I__1213 (
            .O(N__6461),
            .I(N__6455));
    LocalMux I__1212 (
            .O(N__6458),
            .I(\Debounce_SW2.r_CountZ0Z_3 ));
    LocalMux I__1211 (
            .O(N__6455),
            .I(\Debounce_SW2.r_CountZ0Z_3 ));
    InMux I__1210 (
            .O(N__6450),
            .I(N__6445));
    InMux I__1209 (
            .O(N__6449),
            .I(N__6442));
    InMux I__1208 (
            .O(N__6448),
            .I(N__6439));
    LocalMux I__1207 (
            .O(N__6445),
            .I(\Debounce_SW2.r_CountZ0Z_6 ));
    LocalMux I__1206 (
            .O(N__6442),
            .I(\Debounce_SW2.r_CountZ0Z_6 ));
    LocalMux I__1205 (
            .O(N__6439),
            .I(\Debounce_SW2.r_CountZ0Z_6 ));
    CascadeMux I__1204 (
            .O(N__6432),
            .I(\Debounce_SW2.r_Count13_10_cascade_ ));
    InMux I__1203 (
            .O(N__6429),
            .I(N__6424));
    InMux I__1202 (
            .O(N__6428),
            .I(N__6421));
    InMux I__1201 (
            .O(N__6427),
            .I(N__6418));
    LocalMux I__1200 (
            .O(N__6424),
            .I(\Debounce_SW2.r_CountZ0Z_4 ));
    LocalMux I__1199 (
            .O(N__6421),
            .I(\Debounce_SW2.r_CountZ0Z_4 ));
    LocalMux I__1198 (
            .O(N__6418),
            .I(\Debounce_SW2.r_CountZ0Z_4 ));
    InMux I__1197 (
            .O(N__6411),
            .I(N__6407));
    InMux I__1196 (
            .O(N__6410),
            .I(N__6404));
    LocalMux I__1195 (
            .O(N__6407),
            .I(\Debounce_SW2.r_CountZ0Z_11 ));
    LocalMux I__1194 (
            .O(N__6404),
            .I(\Debounce_SW2.r_CountZ0Z_11 ));
    InMux I__1193 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1192 (
            .O(N__6396),
            .I(\Game_Inst.r_Pattern_1_Z0Z_1 ));
    InMux I__1191 (
            .O(N__6393),
            .I(N__6390));
    LocalMux I__1190 (
            .O(N__6390),
            .I(\Game_Inst.r_Pattern_0_Z0Z_0 ));
    InMux I__1189 (
            .O(N__6387),
            .I(N__6384));
    LocalMux I__1188 (
            .O(N__6384),
            .I(\Game_Inst.r_Pattern_1_Z0Z_0 ));
    InMux I__1187 (
            .O(N__6381),
            .I(N__6378));
    LocalMux I__1186 (
            .O(N__6378),
            .I(\Game_Inst.r_Pattern_2_Z0Z_0 ));
    InMux I__1185 (
            .O(N__6375),
            .I(N__6372));
    LocalMux I__1184 (
            .O(N__6372),
            .I(\Game_Inst.r_Pattern_3_Z0Z_0 ));
    InMux I__1183 (
            .O(N__6369),
            .I(N__6365));
    InMux I__1182 (
            .O(N__6368),
            .I(N__6362));
    LocalMux I__1181 (
            .O(N__6365),
            .I(\Game_Inst.w_LFSR_Data_3 ));
    LocalMux I__1180 (
            .O(N__6362),
            .I(\Game_Inst.w_LFSR_Data_3 ));
    InMux I__1179 (
            .O(N__6357),
            .I(N__6354));
    LocalMux I__1178 (
            .O(N__6354),
            .I(\Game_Inst.r_Pattern_6__RNIPJCKZ0Z_1 ));
    InMux I__1177 (
            .O(N__6351),
            .I(N__6347));
    InMux I__1176 (
            .O(N__6350),
            .I(N__6344));
    LocalMux I__1175 (
            .O(N__6347),
            .I(\Game_Inst.w_LFSR_Data_4 ));
    LocalMux I__1174 (
            .O(N__6344),
            .I(\Game_Inst.w_LFSR_Data_4 ));
    InMux I__1173 (
            .O(N__6339),
            .I(N__6336));
    LocalMux I__1172 (
            .O(N__6336),
            .I(\Debounce_SW4.un1_r_Count_8lto11_1 ));
    InMux I__1171 (
            .O(N__6333),
            .I(N__6330));
    LocalMux I__1170 (
            .O(N__6330),
            .I(N__6327));
    Odrv4 I__1169 (
            .O(N__6327),
            .I(\Debounce_SW4.un1_r_Count_8lto17_2 ));
    CascadeMux I__1168 (
            .O(N__6324),
            .I(N__6321));
    InMux I__1167 (
            .O(N__6321),
            .I(N__6318));
    LocalMux I__1166 (
            .O(N__6318),
            .I(\Debounce_SW4.r_Count13_5 ));
    InMux I__1165 (
            .O(N__6315),
            .I(N__6312));
    LocalMux I__1164 (
            .O(N__6312),
            .I(\Debounce_SW4.r_Count13_6 ));
    CascadeMux I__1163 (
            .O(N__6309),
            .I(N__6306));
    InMux I__1162 (
            .O(N__6306),
            .I(N__6303));
    LocalMux I__1161 (
            .O(N__6303),
            .I(\Game_Inst.r_Pattern_1__RNID33IZ0Z_1 ));
    InMux I__1160 (
            .O(N__6300),
            .I(N__6297));
    LocalMux I__1159 (
            .O(N__6297),
            .I(\Game_Inst.r_Pattern_2__RNIHJRIZ0Z_1 ));
    InMux I__1158 (
            .O(N__6294),
            .I(N__6291));
    LocalMux I__1157 (
            .O(N__6291),
            .I(\Game_Inst.r_Pattern_0_Z0Z_1 ));
    InMux I__1156 (
            .O(N__6288),
            .I(N__6285));
    LocalMux I__1155 (
            .O(N__6285),
            .I(\Game_Inst.r_Pattern_2_Z0Z_1 ));
    InMux I__1154 (
            .O(N__6282),
            .I(N__6279));
    LocalMux I__1153 (
            .O(N__6279),
            .I(\Game_Inst.r_Pattern_3_Z0Z_1 ));
    InMux I__1152 (
            .O(N__6276),
            .I(\Debounce_SW2.r_Count_1_cry_15 ));
    InMux I__1151 (
            .O(N__6273),
            .I(bfn_6_15_0_));
    IoInMux I__1150 (
            .O(N__6270),
            .I(N__6267));
    LocalMux I__1149 (
            .O(N__6267),
            .I(N__6264));
    Odrv4 I__1148 (
            .O(N__6264),
            .I(\Debounce_SW4.r_Count12_i ));
    InMux I__1147 (
            .O(N__6261),
            .I(N__6258));
    LocalMux I__1146 (
            .O(N__6258),
            .I(N__6254));
    CascadeMux I__1145 (
            .O(N__6257),
            .I(N__6251));
    Span4Mux_h I__1144 (
            .O(N__6254),
            .I(N__6248));
    InMux I__1143 (
            .O(N__6251),
            .I(N__6245));
    IoSpan4Mux I__1142 (
            .O(N__6248),
            .I(N__6242));
    LocalMux I__1141 (
            .O(N__6245),
            .I(N__6239));
    Odrv4 I__1140 (
            .O(N__6242),
            .I(i_Switch_4_c));
    Odrv12 I__1139 (
            .O(N__6239),
            .I(i_Switch_4_c));
    InMux I__1138 (
            .O(N__6234),
            .I(N__6231));
    LocalMux I__1137 (
            .O(N__6231),
            .I(\Debounce_SW4.r_Count13_10_2 ));
    CascadeMux I__1136 (
            .O(N__6228),
            .I(\Debounce_SW4.r_Count13_9_cascade_ ));
    InMux I__1135 (
            .O(N__6225),
            .I(N__6222));
    LocalMux I__1134 (
            .O(N__6222),
            .I(\Debounce_SW4.r_Count13_1 ));
    CascadeMux I__1133 (
            .O(N__6219),
            .I(\Debounce_SW4.r_Count13_1_cascade_ ));
    CascadeMux I__1132 (
            .O(N__6216),
            .I(\Debounce_SW4.un1_r_Count_8lt11_0_cascade_ ));
    InMux I__1131 (
            .O(N__6213),
            .I(N__6210));
    LocalMux I__1130 (
            .O(N__6210),
            .I(\Debounce_SW4.un1_r_Count_8lt17 ));
    InMux I__1129 (
            .O(N__6207),
            .I(\Debounce_SW2.r_Count_1_cry_6 ));
    InMux I__1128 (
            .O(N__6204),
            .I(\Debounce_SW2.r_Count_1_cry_7 ));
    InMux I__1127 (
            .O(N__6201),
            .I(bfn_6_14_0_));
    InMux I__1126 (
            .O(N__6198),
            .I(\Debounce_SW2.r_Count_1_cry_9 ));
    InMux I__1125 (
            .O(N__6195),
            .I(\Debounce_SW2.r_Count_1_cry_10 ));
    InMux I__1124 (
            .O(N__6192),
            .I(\Debounce_SW2.r_Count_1_cry_11 ));
    InMux I__1123 (
            .O(N__6189),
            .I(\Debounce_SW2.r_Count_1_cry_12 ));
    InMux I__1122 (
            .O(N__6186),
            .I(\Debounce_SW2.r_Count_1_cry_13 ));
    InMux I__1121 (
            .O(N__6183),
            .I(\Debounce_SW2.r_Count_1_cry_14 ));
    InMux I__1120 (
            .O(N__6180),
            .I(N__6177));
    LocalMux I__1119 (
            .O(N__6177),
            .I(\Game_Inst.r_Button_IDZ0Z_0 ));
    InMux I__1118 (
            .O(N__6174),
            .I(N__6169));
    InMux I__1117 (
            .O(N__6173),
            .I(N__6164));
    InMux I__1116 (
            .O(N__6172),
            .I(N__6164));
    LocalMux I__1115 (
            .O(N__6169),
            .I(N__6158));
    LocalMux I__1114 (
            .O(N__6164),
            .I(N__6155));
    InMux I__1113 (
            .O(N__6163),
            .I(N__6152));
    InMux I__1112 (
            .O(N__6162),
            .I(N__6147));
    InMux I__1111 (
            .O(N__6161),
            .I(N__6147));
    Odrv4 I__1110 (
            .O(N__6158),
            .I(\Game_Inst.N_270_li ));
    Odrv4 I__1109 (
            .O(N__6155),
            .I(\Game_Inst.N_270_li ));
    LocalMux I__1108 (
            .O(N__6152),
            .I(\Game_Inst.N_270_li ));
    LocalMux I__1107 (
            .O(N__6147),
            .I(\Game_Inst.N_270_li ));
    CascadeMux I__1106 (
            .O(N__6138),
            .I(N__6135));
    InMux I__1105 (
            .O(N__6135),
            .I(N__6128));
    InMux I__1104 (
            .O(N__6134),
            .I(N__6128));
    CascadeMux I__1103 (
            .O(N__6133),
            .I(N__6125));
    LocalMux I__1102 (
            .O(N__6128),
            .I(N__6122));
    InMux I__1101 (
            .O(N__6125),
            .I(N__6119));
    Odrv12 I__1100 (
            .O(N__6122),
            .I(\Game_Inst.r_SwitchZ0Z_1 ));
    LocalMux I__1099 (
            .O(N__6119),
            .I(\Game_Inst.r_SwitchZ0Z_1 ));
    InMux I__1098 (
            .O(N__6114),
            .I(N__6109));
    InMux I__1097 (
            .O(N__6113),
            .I(N__6104));
    InMux I__1096 (
            .O(N__6112),
            .I(N__6100));
    LocalMux I__1095 (
            .O(N__6109),
            .I(N__6097));
    InMux I__1094 (
            .O(N__6108),
            .I(N__6094));
    InMux I__1093 (
            .O(N__6107),
            .I(N__6091));
    LocalMux I__1092 (
            .O(N__6104),
            .I(N__6083));
    CascadeMux I__1091 (
            .O(N__6103),
            .I(N__6080));
    LocalMux I__1090 (
            .O(N__6100),
            .I(N__6077));
    Span4Mux_v I__1089 (
            .O(N__6097),
            .I(N__6070));
    LocalMux I__1088 (
            .O(N__6094),
            .I(N__6070));
    LocalMux I__1087 (
            .O(N__6091),
            .I(N__6070));
    InMux I__1086 (
            .O(N__6090),
            .I(N__6067));
    InMux I__1085 (
            .O(N__6089),
            .I(N__6060));
    InMux I__1084 (
            .O(N__6088),
            .I(N__6060));
    InMux I__1083 (
            .O(N__6087),
            .I(N__6060));
    InMux I__1082 (
            .O(N__6086),
            .I(N__6057));
    Span4Mux_h I__1081 (
            .O(N__6083),
            .I(N__6054));
    InMux I__1080 (
            .O(N__6080),
            .I(N__6051));
    Span4Mux_h I__1079 (
            .O(N__6077),
            .I(N__6048));
    Span4Mux_h I__1078 (
            .O(N__6070),
            .I(N__6045));
    LocalMux I__1077 (
            .O(N__6067),
            .I(N__6040));
    LocalMux I__1076 (
            .O(N__6060),
            .I(N__6040));
    LocalMux I__1075 (
            .O(N__6057),
            .I(w_Switch_1));
    Odrv4 I__1074 (
            .O(N__6054),
            .I(w_Switch_1));
    LocalMux I__1073 (
            .O(N__6051),
            .I(w_Switch_1));
    Odrv4 I__1072 (
            .O(N__6048),
            .I(w_Switch_1));
    Odrv4 I__1071 (
            .O(N__6045),
            .I(w_Switch_1));
    Odrv12 I__1070 (
            .O(N__6040),
            .I(w_Switch_1));
    InMux I__1069 (
            .O(N__6027),
            .I(N__6024));
    LocalMux I__1068 (
            .O(N__6024),
            .I(N__6021));
    Odrv4 I__1067 (
            .O(N__6021),
            .I(\Game_Inst.r_Button_IDZ0Z_1 ));
    InMux I__1066 (
            .O(N__6018),
            .I(\Debounce_SW2.r_Count_1_cry_1 ));
    InMux I__1065 (
            .O(N__6015),
            .I(\Debounce_SW2.r_Count_1_cry_2 ));
    InMux I__1064 (
            .O(N__6012),
            .I(\Debounce_SW2.r_Count_1_cry_3 ));
    InMux I__1063 (
            .O(N__6009),
            .I(\Debounce_SW2.r_Count_1_cry_4 ));
    InMux I__1062 (
            .O(N__6006),
            .I(\Debounce_SW2.r_Count_1_cry_5 ));
    InMux I__1061 (
            .O(N__6003),
            .I(N__5996));
    InMux I__1060 (
            .O(N__6002),
            .I(N__5993));
    InMux I__1059 (
            .O(N__6001),
            .I(N__5990));
    InMux I__1058 (
            .O(N__6000),
            .I(N__5985));
    InMux I__1057 (
            .O(N__5999),
            .I(N__5985));
    LocalMux I__1056 (
            .O(N__5996),
            .I(\Game_Inst.r_IndexZ1Z_1 ));
    LocalMux I__1055 (
            .O(N__5993),
            .I(\Game_Inst.r_IndexZ1Z_1 ));
    LocalMux I__1054 (
            .O(N__5990),
            .I(\Game_Inst.r_IndexZ1Z_1 ));
    LocalMux I__1053 (
            .O(N__5985),
            .I(\Game_Inst.r_IndexZ1Z_1 ));
    InMux I__1052 (
            .O(N__5976),
            .I(N__5972));
    InMux I__1051 (
            .O(N__5975),
            .I(N__5969));
    LocalMux I__1050 (
            .O(N__5972),
            .I(N__5966));
    LocalMux I__1049 (
            .O(N__5969),
            .I(\Game_Inst.N_276_0 ));
    Odrv4 I__1048 (
            .O(N__5966),
            .I(\Game_Inst.N_276_0 ));
    InMux I__1047 (
            .O(N__5961),
            .I(N__5953));
    InMux I__1046 (
            .O(N__5960),
            .I(N__5948));
    InMux I__1045 (
            .O(N__5959),
            .I(N__5948));
    InMux I__1044 (
            .O(N__5958),
            .I(N__5941));
    InMux I__1043 (
            .O(N__5957),
            .I(N__5941));
    InMux I__1042 (
            .O(N__5956),
            .I(N__5941));
    LocalMux I__1041 (
            .O(N__5953),
            .I(\Game_Inst.r_IndexZ0Z_2 ));
    LocalMux I__1040 (
            .O(N__5948),
            .I(\Game_Inst.r_IndexZ0Z_2 ));
    LocalMux I__1039 (
            .O(N__5941),
            .I(\Game_Inst.r_IndexZ0Z_2 ));
    CascadeMux I__1038 (
            .O(N__5934),
            .I(\Game_Inst.r_Pattern_5__RNIL3KJZ0Z_1_cascade_ ));
    InMux I__1037 (
            .O(N__5931),
            .I(N__5928));
    LocalMux I__1036 (
            .O(N__5928),
            .I(\Game_Inst.un1_r_Pattern_0__7_ns_1_1 ));
    CascadeMux I__1035 (
            .O(N__5925),
            .I(\Game_Inst.N_31_cascade_ ));
    InMux I__1034 (
            .O(N__5922),
            .I(N__5916));
    InMux I__1033 (
            .O(N__5921),
            .I(N__5916));
    LocalMux I__1032 (
            .O(N__5916),
            .I(N__5911));
    InMux I__1031 (
            .O(N__5915),
            .I(N__5908));
    InMux I__1030 (
            .O(N__5914),
            .I(N__5905));
    Odrv4 I__1029 (
            .O(N__5911),
            .I(\Game_Inst.un1_r_Pattern_0__1_i_0 ));
    LocalMux I__1028 (
            .O(N__5908),
            .I(\Game_Inst.un1_r_Pattern_0__1_i_0 ));
    LocalMux I__1027 (
            .O(N__5905),
            .I(\Game_Inst.un1_r_Pattern_0__1_i_0 ));
    CascadeMux I__1026 (
            .O(N__5898),
            .I(N__5895));
    InMux I__1025 (
            .O(N__5895),
            .I(N__5889));
    InMux I__1024 (
            .O(N__5894),
            .I(N__5889));
    LocalMux I__1023 (
            .O(N__5889),
            .I(\Game_Inst.N_311 ));
    InMux I__1022 (
            .O(N__5886),
            .I(N__5880));
    CascadeMux I__1021 (
            .O(N__5885),
            .I(N__5877));
    CascadeMux I__1020 (
            .O(N__5884),
            .I(N__5873));
    CascadeMux I__1019 (
            .O(N__5883),
            .I(N__5862));
    LocalMux I__1018 (
            .O(N__5880),
            .I(N__5859));
    InMux I__1017 (
            .O(N__5877),
            .I(N__5854));
    InMux I__1016 (
            .O(N__5876),
            .I(N__5854));
    InMux I__1015 (
            .O(N__5873),
            .I(N__5851));
    InMux I__1014 (
            .O(N__5872),
            .I(N__5846));
    InMux I__1013 (
            .O(N__5871),
            .I(N__5846));
    InMux I__1012 (
            .O(N__5870),
            .I(N__5843));
    InMux I__1011 (
            .O(N__5869),
            .I(N__5838));
    InMux I__1010 (
            .O(N__5868),
            .I(N__5838));
    InMux I__1009 (
            .O(N__5867),
            .I(N__5835));
    InMux I__1008 (
            .O(N__5866),
            .I(N__5829));
    InMux I__1007 (
            .O(N__5865),
            .I(N__5829));
    InMux I__1006 (
            .O(N__5862),
            .I(N__5826));
    Span4Mux_v I__1005 (
            .O(N__5859),
            .I(N__5817));
    LocalMux I__1004 (
            .O(N__5854),
            .I(N__5817));
    LocalMux I__1003 (
            .O(N__5851),
            .I(N__5817));
    LocalMux I__1002 (
            .O(N__5846),
            .I(N__5817));
    LocalMux I__1001 (
            .O(N__5843),
            .I(N__5812));
    LocalMux I__1000 (
            .O(N__5838),
            .I(N__5812));
    LocalMux I__999 (
            .O(N__5835),
            .I(N__5809));
    InMux I__998 (
            .O(N__5834),
            .I(N__5806));
    LocalMux I__997 (
            .O(N__5829),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    LocalMux I__996 (
            .O(N__5826),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    Odrv4 I__995 (
            .O(N__5817),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    Odrv12 I__994 (
            .O(N__5812),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    Odrv4 I__993 (
            .O(N__5809),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    LocalMux I__992 (
            .O(N__5806),
            .I(\Game_Inst.r_SM_MainZ0Z_2 ));
    CascadeMux I__991 (
            .O(N__5793),
            .I(\Game_Inst.un1_r_Pattern_0__1_i_0_cascade_ ));
    InMux I__990 (
            .O(N__5790),
            .I(N__5783));
    InMux I__989 (
            .O(N__5789),
            .I(N__5783));
    InMux I__988 (
            .O(N__5788),
            .I(N__5780));
    LocalMux I__987 (
            .O(N__5783),
            .I(N__5777));
    LocalMux I__986 (
            .O(N__5780),
            .I(N__5772));
    Span4Mux_h I__985 (
            .O(N__5777),
            .I(N__5772));
    Odrv4 I__984 (
            .O(N__5772),
            .I(\Game_Inst.N_309 ));
    InMux I__983 (
            .O(N__5769),
            .I(N__5759));
    InMux I__982 (
            .O(N__5768),
            .I(N__5759));
    InMux I__981 (
            .O(N__5767),
            .I(N__5756));
    InMux I__980 (
            .O(N__5766),
            .I(N__5751));
    InMux I__979 (
            .O(N__5765),
            .I(N__5751));
    InMux I__978 (
            .O(N__5764),
            .I(N__5742));
    LocalMux I__977 (
            .O(N__5759),
            .I(N__5739));
    LocalMux I__976 (
            .O(N__5756),
            .I(N__5734));
    LocalMux I__975 (
            .O(N__5751),
            .I(N__5734));
    InMux I__974 (
            .O(N__5750),
            .I(N__5731));
    InMux I__973 (
            .O(N__5749),
            .I(N__5728));
    InMux I__972 (
            .O(N__5748),
            .I(N__5719));
    InMux I__971 (
            .O(N__5747),
            .I(N__5719));
    InMux I__970 (
            .O(N__5746),
            .I(N__5719));
    InMux I__969 (
            .O(N__5745),
            .I(N__5719));
    LocalMux I__968 (
            .O(N__5742),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    Odrv4 I__967 (
            .O(N__5739),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    Odrv4 I__966 (
            .O(N__5734),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    LocalMux I__965 (
            .O(N__5731),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    LocalMux I__964 (
            .O(N__5728),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    LocalMux I__963 (
            .O(N__5719),
            .I(\Game_Inst.r_SM_MainZ0Z_1 ));
    CascadeMux I__962 (
            .O(N__5706),
            .I(\Game_Inst.N_269_0_cascade_ ));
    InMux I__961 (
            .O(N__5703),
            .I(N__5698));
    InMux I__960 (
            .O(N__5702),
            .I(N__5693));
    InMux I__959 (
            .O(N__5701),
            .I(N__5693));
    LocalMux I__958 (
            .O(N__5698),
            .I(\Game_Inst.N_314 ));
    LocalMux I__957 (
            .O(N__5693),
            .I(\Game_Inst.N_314 ));
    InMux I__956 (
            .O(N__5688),
            .I(N__5685));
    LocalMux I__955 (
            .O(N__5685),
            .I(\Game_Inst.r_SwitchZ0Z_4 ));
    InMux I__954 (
            .O(N__5682),
            .I(N__5678));
    InMux I__953 (
            .O(N__5681),
            .I(N__5673));
    LocalMux I__952 (
            .O(N__5678),
            .I(N__5670));
    InMux I__951 (
            .O(N__5677),
            .I(N__5667));
    InMux I__950 (
            .O(N__5676),
            .I(N__5664));
    LocalMux I__949 (
            .O(N__5673),
            .I(N__5651));
    Span4Mux_h I__948 (
            .O(N__5670),
            .I(N__5648));
    LocalMux I__947 (
            .O(N__5667),
            .I(N__5643));
    LocalMux I__946 (
            .O(N__5664),
            .I(N__5643));
    InMux I__945 (
            .O(N__5663),
            .I(N__5638));
    InMux I__944 (
            .O(N__5662),
            .I(N__5638));
    InMux I__943 (
            .O(N__5661),
            .I(N__5635));
    InMux I__942 (
            .O(N__5660),
            .I(N__5628));
    InMux I__941 (
            .O(N__5659),
            .I(N__5628));
    InMux I__940 (
            .O(N__5658),
            .I(N__5628));
    InMux I__939 (
            .O(N__5657),
            .I(N__5619));
    InMux I__938 (
            .O(N__5656),
            .I(N__5619));
    InMux I__937 (
            .O(N__5655),
            .I(N__5619));
    InMux I__936 (
            .O(N__5654),
            .I(N__5619));
    Odrv4 I__935 (
            .O(N__5651),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    Odrv4 I__934 (
            .O(N__5648),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    Odrv4 I__933 (
            .O(N__5643),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    LocalMux I__932 (
            .O(N__5638),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    LocalMux I__931 (
            .O(N__5635),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    LocalMux I__930 (
            .O(N__5628),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    LocalMux I__929 (
            .O(N__5619),
            .I(\Game_Inst.r_SM_MainZ0Z_0 ));
    InMux I__928 (
            .O(N__5604),
            .I(N__5600));
    InMux I__927 (
            .O(N__5603),
            .I(N__5597));
    LocalMux I__926 (
            .O(N__5600),
            .I(\Game_Inst.N_275_0 ));
    LocalMux I__925 (
            .O(N__5597),
            .I(\Game_Inst.N_275_0 ));
    CascadeMux I__924 (
            .O(N__5592),
            .I(\Game_Inst.N_275_0_cascade_ ));
    CascadeMux I__923 (
            .O(N__5589),
            .I(\Game_Inst.N_268_0_cascade_ ));
    InMux I__922 (
            .O(N__5586),
            .I(N__5581));
    InMux I__921 (
            .O(N__5585),
            .I(N__5576));
    InMux I__920 (
            .O(N__5584),
            .I(N__5576));
    LocalMux I__919 (
            .O(N__5581),
            .I(\Game_Inst.r_Index_0_sqmuxa ));
    LocalMux I__918 (
            .O(N__5576),
            .I(\Game_Inst.r_Index_0_sqmuxa ));
    CascadeMux I__917 (
            .O(N__5571),
            .I(\Game_Inst.r_Pattern_1__RNIB13IZ0Z_0_cascade_ ));
    InMux I__916 (
            .O(N__5568),
            .I(N__5565));
    LocalMux I__915 (
            .O(N__5565),
            .I(\Game_Inst.r_Pattern_2__RNIFHRIZ0Z_0 ));
    InMux I__914 (
            .O(N__5562),
            .I(N__5559));
    LocalMux I__913 (
            .O(N__5559),
            .I(\Game_Inst.SUM_i_o3_1_0 ));
    InMux I__912 (
            .O(N__5556),
            .I(N__5553));
    LocalMux I__911 (
            .O(N__5553),
            .I(\Game_Inst.un1_r_Pattern_0__7_ns_1_0 ));
    CascadeMux I__910 (
            .O(N__5550),
            .I(\Game_Inst.N_287_0_cascade_ ));
    InMux I__909 (
            .O(N__5547),
            .I(N__5541));
    InMux I__908 (
            .O(N__5546),
            .I(N__5541));
    LocalMux I__907 (
            .O(N__5541),
            .I(\Game_Inst.N_262_0 ));
    InMux I__906 (
            .O(N__5538),
            .I(N__5535));
    LocalMux I__905 (
            .O(N__5535),
            .I(\Game_Inst.o_Score_RNO_0Z0Z_1 ));
    CascadeMux I__904 (
            .O(N__5532),
            .I(N__5526));
    InMux I__903 (
            .O(N__5531),
            .I(N__5521));
    InMux I__902 (
            .O(N__5530),
            .I(N__5521));
    InMux I__901 (
            .O(N__5529),
            .I(N__5516));
    InMux I__900 (
            .O(N__5526),
            .I(N__5516));
    LocalMux I__899 (
            .O(N__5521),
            .I(\Game_Inst.N_287_0 ));
    LocalMux I__898 (
            .O(N__5516),
            .I(\Game_Inst.N_287_0 ));
    CascadeMux I__897 (
            .O(N__5511),
            .I(N__5505));
    InMux I__896 (
            .O(N__5510),
            .I(N__5501));
    InMux I__895 (
            .O(N__5509),
            .I(N__5498));
    InMux I__894 (
            .O(N__5508),
            .I(N__5493));
    InMux I__893 (
            .O(N__5505),
            .I(N__5493));
    InMux I__892 (
            .O(N__5504),
            .I(N__5490));
    LocalMux I__891 (
            .O(N__5501),
            .I(\Game_Inst.o_Score_0_sqmuxa ));
    LocalMux I__890 (
            .O(N__5498),
            .I(\Game_Inst.o_Score_0_sqmuxa ));
    LocalMux I__889 (
            .O(N__5493),
            .I(\Game_Inst.o_Score_0_sqmuxa ));
    LocalMux I__888 (
            .O(N__5490),
            .I(\Game_Inst.o_Score_0_sqmuxa ));
    InMux I__887 (
            .O(N__5481),
            .I(N__5475));
    InMux I__886 (
            .O(N__5480),
            .I(N__5475));
    LocalMux I__885 (
            .O(N__5475),
            .I(N__5470));
    InMux I__884 (
            .O(N__5474),
            .I(N__5467));
    InMux I__883 (
            .O(N__5473),
            .I(N__5464));
    Odrv4 I__882 (
            .O(N__5470),
            .I(\Game_Inst.N_310 ));
    LocalMux I__881 (
            .O(N__5467),
            .I(\Game_Inst.N_310 ));
    LocalMux I__880 (
            .O(N__5464),
            .I(\Game_Inst.N_310 ));
    InMux I__879 (
            .O(N__5457),
            .I(N__5443));
    InMux I__878 (
            .O(N__5456),
            .I(N__5443));
    InMux I__877 (
            .O(N__5455),
            .I(N__5443));
    InMux I__876 (
            .O(N__5454),
            .I(N__5443));
    InMux I__875 (
            .O(N__5453),
            .I(N__5440));
    InMux I__874 (
            .O(N__5452),
            .I(N__5436));
    LocalMux I__873 (
            .O(N__5443),
            .I(N__5433));
    LocalMux I__872 (
            .O(N__5440),
            .I(N__5430));
    InMux I__871 (
            .O(N__5439),
            .I(N__5427));
    LocalMux I__870 (
            .O(N__5436),
            .I(N__5421));
    Span4Mux_s3_v I__869 (
            .O(N__5433),
            .I(N__5414));
    Span4Mux_s3_v I__868 (
            .O(N__5430),
            .I(N__5414));
    LocalMux I__867 (
            .O(N__5427),
            .I(N__5414));
    InMux I__866 (
            .O(N__5426),
            .I(N__5411));
    InMux I__865 (
            .O(N__5425),
            .I(N__5408));
    InMux I__864 (
            .O(N__5424),
            .I(N__5405));
    Odrv12 I__863 (
            .O(N__5421),
            .I(w_Score_1));
    Odrv4 I__862 (
            .O(N__5414),
            .I(w_Score_1));
    LocalMux I__861 (
            .O(N__5411),
            .I(w_Score_1));
    LocalMux I__860 (
            .O(N__5408),
            .I(w_Score_1));
    LocalMux I__859 (
            .O(N__5405),
            .I(w_Score_1));
    CascadeMux I__858 (
            .O(N__5394),
            .I(N__5386));
    CascadeMux I__857 (
            .O(N__5393),
            .I(N__5383));
    CascadeMux I__856 (
            .O(N__5392),
            .I(N__5380));
    InMux I__855 (
            .O(N__5391),
            .I(N__5376));
    InMux I__854 (
            .O(N__5390),
            .I(N__5373));
    InMux I__853 (
            .O(N__5389),
            .I(N__5363));
    InMux I__852 (
            .O(N__5386),
            .I(N__5363));
    InMux I__851 (
            .O(N__5383),
            .I(N__5363));
    InMux I__850 (
            .O(N__5380),
            .I(N__5363));
    InMux I__849 (
            .O(N__5379),
            .I(N__5360));
    LocalMux I__848 (
            .O(N__5376),
            .I(N__5355));
    LocalMux I__847 (
            .O(N__5373),
            .I(N__5355));
    CascadeMux I__846 (
            .O(N__5372),
            .I(N__5351));
    LocalMux I__845 (
            .O(N__5363),
            .I(N__5347));
    LocalMux I__844 (
            .O(N__5360),
            .I(N__5342));
    Span4Mux_s3_v I__843 (
            .O(N__5355),
            .I(N__5342));
    InMux I__842 (
            .O(N__5354),
            .I(N__5339));
    InMux I__841 (
            .O(N__5351),
            .I(N__5336));
    InMux I__840 (
            .O(N__5350),
            .I(N__5333));
    Odrv12 I__839 (
            .O(N__5347),
            .I(w_Score_2));
    Odrv4 I__838 (
            .O(N__5342),
            .I(w_Score_2));
    LocalMux I__837 (
            .O(N__5339),
            .I(w_Score_2));
    LocalMux I__836 (
            .O(N__5336),
            .I(w_Score_2));
    LocalMux I__835 (
            .O(N__5333),
            .I(w_Score_2));
    CascadeMux I__834 (
            .O(N__5322),
            .I(N__5313));
    CascadeMux I__833 (
            .O(N__5321),
            .I(N__5310));
    CascadeMux I__832 (
            .O(N__5320),
            .I(N__5307));
    CascadeMux I__831 (
            .O(N__5319),
            .I(N__5304));
    InMux I__830 (
            .O(N__5318),
            .I(N__5295));
    InMux I__829 (
            .O(N__5317),
            .I(N__5295));
    InMux I__828 (
            .O(N__5316),
            .I(N__5295));
    InMux I__827 (
            .O(N__5313),
            .I(N__5295));
    InMux I__826 (
            .O(N__5310),
            .I(N__5292));
    InMux I__825 (
            .O(N__5307),
            .I(N__5289));
    InMux I__824 (
            .O(N__5304),
            .I(N__5283));
    LocalMux I__823 (
            .O(N__5295),
            .I(N__5276));
    LocalMux I__822 (
            .O(N__5292),
            .I(N__5276));
    LocalMux I__821 (
            .O(N__5289),
            .I(N__5276));
    InMux I__820 (
            .O(N__5288),
            .I(N__5273));
    CascadeMux I__819 (
            .O(N__5287),
            .I(N__5270));
    InMux I__818 (
            .O(N__5286),
            .I(N__5267));
    LocalMux I__817 (
            .O(N__5283),
            .I(N__5260));
    Span4Mux_v I__816 (
            .O(N__5276),
            .I(N__5260));
    LocalMux I__815 (
            .O(N__5273),
            .I(N__5260));
    InMux I__814 (
            .O(N__5270),
            .I(N__5257));
    LocalMux I__813 (
            .O(N__5267),
            .I(w_Score_3));
    Odrv4 I__812 (
            .O(N__5260),
            .I(w_Score_3));
    LocalMux I__811 (
            .O(N__5257),
            .I(w_Score_3));
    InMux I__810 (
            .O(N__5250),
            .I(N__5247));
    LocalMux I__809 (
            .O(N__5247),
            .I(N__5238));
    InMux I__808 (
            .O(N__5246),
            .I(N__5229));
    InMux I__807 (
            .O(N__5245),
            .I(N__5229));
    InMux I__806 (
            .O(N__5244),
            .I(N__5229));
    InMux I__805 (
            .O(N__5243),
            .I(N__5229));
    InMux I__804 (
            .O(N__5242),
            .I(N__5226));
    InMux I__803 (
            .O(N__5241),
            .I(N__5223));
    Span4Mux_v I__802 (
            .O(N__5238),
            .I(N__5217));
    LocalMux I__801 (
            .O(N__5229),
            .I(N__5212));
    LocalMux I__800 (
            .O(N__5226),
            .I(N__5212));
    LocalMux I__799 (
            .O(N__5223),
            .I(N__5209));
    InMux I__798 (
            .O(N__5222),
            .I(N__5206));
    InMux I__797 (
            .O(N__5221),
            .I(N__5203));
    InMux I__796 (
            .O(N__5220),
            .I(N__5200));
    Odrv4 I__795 (
            .O(N__5217),
            .I(w_Score_0));
    Odrv12 I__794 (
            .O(N__5212),
            .I(w_Score_0));
    Odrv4 I__793 (
            .O(N__5209),
            .I(w_Score_0));
    LocalMux I__792 (
            .O(N__5206),
            .I(w_Score_0));
    LocalMux I__791 (
            .O(N__5203),
            .I(w_Score_0));
    LocalMux I__790 (
            .O(N__5200),
            .I(w_Score_0));
    IoInMux I__789 (
            .O(N__5187),
            .I(N__5184));
    LocalMux I__788 (
            .O(N__5184),
            .I(r_Hex_Encoding_i_2));
    CascadeMux I__787 (
            .O(N__5181),
            .I(N__5177));
    InMux I__786 (
            .O(N__5180),
            .I(N__5174));
    InMux I__785 (
            .O(N__5177),
            .I(N__5170));
    LocalMux I__784 (
            .O(N__5174),
            .I(N__5166));
    InMux I__783 (
            .O(N__5173),
            .I(N__5163));
    LocalMux I__782 (
            .O(N__5170),
            .I(N__5160));
    InMux I__781 (
            .O(N__5169),
            .I(N__5157));
    Odrv4 I__780 (
            .O(N__5166),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ));
    LocalMux I__779 (
            .O(N__5163),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ));
    Odrv4 I__778 (
            .O(N__5160),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ));
    LocalMux I__777 (
            .O(N__5157),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ));
    InMux I__776 (
            .O(N__5148),
            .I(N__5143));
    InMux I__775 (
            .O(N__5147),
            .I(N__5140));
    InMux I__774 (
            .O(N__5146),
            .I(N__5137));
    LocalMux I__773 (
            .O(N__5143),
            .I(N__5134));
    LocalMux I__772 (
            .O(N__5140),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_1 ));
    LocalMux I__771 (
            .O(N__5137),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_1 ));
    Odrv4 I__770 (
            .O(N__5134),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_1 ));
    SRMux I__769 (
            .O(N__5127),
            .I(N__5121));
    SRMux I__768 (
            .O(N__5126),
            .I(N__5118));
    SRMux I__767 (
            .O(N__5125),
            .I(N__5115));
    SRMux I__766 (
            .O(N__5124),
            .I(N__5112));
    LocalMux I__765 (
            .O(N__5121),
            .I(N__5109));
    LocalMux I__764 (
            .O(N__5118),
            .I(N__5106));
    LocalMux I__763 (
            .O(N__5115),
            .I(N__5103));
    LocalMux I__762 (
            .O(N__5112),
            .I(N__5100));
    Glb2LocalMux I__761 (
            .O(N__5109),
            .I(N__5091));
    Glb2LocalMux I__760 (
            .O(N__5106),
            .I(N__5091));
    Glb2LocalMux I__759 (
            .O(N__5103),
            .I(N__5091));
    Glb2LocalMux I__758 (
            .O(N__5100),
            .I(N__5091));
    GlobalMux I__757 (
            .O(N__5091),
            .I(N__5088));
    gio2CtrlBuf I__756 (
            .O(N__5088),
            .I(\Game_Inst.Count_Inst.N_213_g ));
    CascadeMux I__755 (
            .O(N__5085),
            .I(\Game_Inst.r_SM_Main_100_d_cascade_ ));
    IoInMux I__754 (
            .O(N__5082),
            .I(N__5079));
    LocalMux I__753 (
            .O(N__5079),
            .I(N__5076));
    Span4Mux_s2_h I__752 (
            .O(N__5076),
            .I(N__5073));
    Span4Mux_h I__751 (
            .O(N__5073),
            .I(N__5070));
    Odrv4 I__750 (
            .O(N__5070),
            .I(Game_Inst_o_LED_1_0_i));
    InMux I__749 (
            .O(N__5067),
            .I(N__5063));
    CascadeMux I__748 (
            .O(N__5066),
            .I(N__5060));
    LocalMux I__747 (
            .O(N__5063),
            .I(N__5057));
    InMux I__746 (
            .O(N__5060),
            .I(N__5054));
    Span4Mux_h I__745 (
            .O(N__5057),
            .I(N__5051));
    LocalMux I__744 (
            .O(N__5054),
            .I(\Game_Inst.N_334_0 ));
    Odrv4 I__743 (
            .O(N__5051),
            .I(\Game_Inst.N_334_0 ));
    CascadeMux I__742 (
            .O(N__5046),
            .I(N__5042));
    InMux I__741 (
            .O(N__5045),
            .I(N__5039));
    InMux I__740 (
            .O(N__5042),
            .I(N__5036));
    LocalMux I__739 (
            .O(N__5039),
            .I(\Game_Inst.r_SM_Main_0_sqmuxa_2_1 ));
    LocalMux I__738 (
            .O(N__5036),
            .I(\Game_Inst.r_SM_Main_0_sqmuxa_2_1 ));
    InMux I__737 (
            .O(N__5031),
            .I(N__5027));
    InMux I__736 (
            .O(N__5030),
            .I(N__5024));
    LocalMux I__735 (
            .O(N__5027),
            .I(\Game_Inst.N_335_0 ));
    LocalMux I__734 (
            .O(N__5024),
            .I(\Game_Inst.N_335_0 ));
    InMux I__733 (
            .O(N__5019),
            .I(N__5016));
    LocalMux I__732 (
            .O(N__5016),
            .I(\Game_Inst.r_SM_Main_ns_i_0_2 ));
    CascadeMux I__731 (
            .O(N__5013),
            .I(\Game_Inst.r_Index16_NE_1_cascade_ ));
    InMux I__730 (
            .O(N__5010),
            .I(N__5001));
    InMux I__729 (
            .O(N__5009),
            .I(N__5001));
    InMux I__728 (
            .O(N__5008),
            .I(N__5001));
    LocalMux I__727 (
            .O(N__5001),
            .I(N__4997));
    InMux I__726 (
            .O(N__5000),
            .I(N__4994));
    Odrv4 I__725 (
            .O(N__4997),
            .I(\Game_Inst.N_330_li ));
    LocalMux I__724 (
            .O(N__4994),
            .I(\Game_Inst.N_330_li ));
    CascadeMux I__723 (
            .O(N__4989),
            .I(\Game_Inst.N_330_li_cascade_ ));
    InMux I__722 (
            .O(N__4986),
            .I(N__4983));
    LocalMux I__721 (
            .O(N__4983),
            .I(N__4980));
    Odrv4 I__720 (
            .O(N__4980),
            .I(\Game_Inst.r_SM_Main_0_sqmuxa_1 ));
    InMux I__719 (
            .O(N__4977),
            .I(N__4971));
    InMux I__718 (
            .O(N__4976),
            .I(N__4968));
    InMux I__717 (
            .O(N__4975),
            .I(N__4965));
    InMux I__716 (
            .O(N__4974),
            .I(N__4962));
    LocalMux I__715 (
            .O(N__4971),
            .I(\Game_Inst.r_Button_DVZ0 ));
    LocalMux I__714 (
            .O(N__4968),
            .I(\Game_Inst.r_Button_DVZ0 ));
    LocalMux I__713 (
            .O(N__4965),
            .I(\Game_Inst.r_Button_DVZ0 ));
    LocalMux I__712 (
            .O(N__4962),
            .I(\Game_Inst.r_Button_DVZ0 ));
    CascadeMux I__711 (
            .O(N__4953),
            .I(\Game_Inst.r_SM_Main_98_d_cascade_ ));
    InMux I__710 (
            .O(N__4950),
            .I(N__4947));
    LocalMux I__709 (
            .O(N__4947),
            .I(\Game_Inst.o_Score_RNO_0Z0Z_0 ));
    InMux I__708 (
            .O(N__4944),
            .I(\Game_Inst.un1_o_Score_cry_0 ));
    InMux I__707 (
            .O(N__4941),
            .I(N__4938));
    LocalMux I__706 (
            .O(N__4938),
            .I(\Game_Inst.o_Score_RNO_0Z0Z_2 ));
    InMux I__705 (
            .O(N__4935),
            .I(\Game_Inst.un1_o_Score_cry_1 ));
    InMux I__704 (
            .O(N__4932),
            .I(\Game_Inst.un1_o_Score_cry_2 ));
    CascadeMux I__703 (
            .O(N__4929),
            .I(\Game_Inst.o_Score_RNO_0Z0Z_3_cascade_ ));
    InMux I__702 (
            .O(N__4926),
            .I(N__4919));
    InMux I__701 (
            .O(N__4925),
            .I(N__4916));
    InMux I__700 (
            .O(N__4924),
            .I(N__4909));
    InMux I__699 (
            .O(N__4923),
            .I(N__4909));
    InMux I__698 (
            .O(N__4922),
            .I(N__4909));
    LocalMux I__697 (
            .O(N__4919),
            .I(\Game_Inst.w_Toggle ));
    LocalMux I__696 (
            .O(N__4916),
            .I(\Game_Inst.w_Toggle ));
    LocalMux I__695 (
            .O(N__4909),
            .I(\Game_Inst.w_Toggle ));
    InMux I__694 (
            .O(N__4902),
            .I(N__4897));
    InMux I__693 (
            .O(N__4901),
            .I(N__4892));
    InMux I__692 (
            .O(N__4900),
            .I(N__4892));
    LocalMux I__691 (
            .O(N__4897),
            .I(\Game_Inst.r_ToggleZ0 ));
    LocalMux I__690 (
            .O(N__4892),
            .I(\Game_Inst.r_ToggleZ0 ));
    InMux I__689 (
            .O(N__4887),
            .I(N__4880));
    InMux I__688 (
            .O(N__4886),
            .I(N__4880));
    InMux I__687 (
            .O(N__4885),
            .I(N__4877));
    LocalMux I__686 (
            .O(N__4880),
            .I(N__4874));
    LocalMux I__685 (
            .O(N__4877),
            .I(\Game_Inst.r_SM_Main7 ));
    Odrv4 I__684 (
            .O(N__4874),
            .I(\Game_Inst.r_SM_Main7 ));
    CascadeMux I__683 (
            .O(N__4869),
            .I(\Game_Inst.r_SM_Main_0_sqmuxa_2_1_cascade_ ));
    InMux I__682 (
            .O(N__4866),
            .I(N__4863));
    LocalMux I__681 (
            .O(N__4863),
            .I(\Game_Inst.N_345 ));
    CascadeMux I__680 (
            .O(N__4860),
            .I(\Game_Inst.N_345_cascade_ ));
    CascadeMux I__679 (
            .O(N__4857),
            .I(\Game_Inst.SUM_i_0_1_cascade_ ));
    InMux I__678 (
            .O(N__4854),
            .I(N__4850));
    InMux I__677 (
            .O(N__4853),
            .I(N__4847));
    LocalMux I__676 (
            .O(N__4850),
            .I(N__4844));
    LocalMux I__675 (
            .O(N__4847),
            .I(N__4841));
    Odrv4 I__674 (
            .O(N__4844),
            .I(\Game_Inst.N_333_0 ));
    Odrv4 I__673 (
            .O(N__4841),
            .I(\Game_Inst.N_333_0 ));
    InMux I__672 (
            .O(N__4836),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_22 ));
    CascadeMux I__671 (
            .O(N__4833),
            .I(N__4829));
    InMux I__670 (
            .O(N__4832),
            .I(N__4826));
    InMux I__669 (
            .O(N__4829),
            .I(N__4823));
    LocalMux I__668 (
            .O(N__4826),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_23 ));
    LocalMux I__667 (
            .O(N__4823),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_23 ));
    CascadeMux I__666 (
            .O(N__4818),
            .I(N__4814));
    InMux I__665 (
            .O(N__4817),
            .I(N__4811));
    InMux I__664 (
            .O(N__4814),
            .I(N__4808));
    LocalMux I__663 (
            .O(N__4811),
            .I(\Game_Inst.r_SM_Main_ns_i_a4_0_0 ));
    LocalMux I__662 (
            .O(N__4808),
            .I(\Game_Inst.r_SM_Main_ns_i_a4_0_0 ));
    CascadeMux I__661 (
            .O(N__4803),
            .I(\Game_Inst.r_SM_Main_ns_i_0_1_cascade_ ));
    CascadeMux I__660 (
            .O(N__4800),
            .I(\Game_Inst.r_SM_Main_ns_i_2_1_cascade_ ));
    InMux I__659 (
            .O(N__4797),
            .I(N__4794));
    LocalMux I__658 (
            .O(N__4794),
            .I(\Game_Inst.r_SM_Main_ns_i_a4_0_1_1 ));
    CascadeMux I__657 (
            .O(N__4791),
            .I(N__4787));
    InMux I__656 (
            .O(N__4790),
            .I(N__4784));
    InMux I__655 (
            .O(N__4787),
            .I(N__4781));
    LocalMux I__654 (
            .O(N__4784),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_14 ));
    LocalMux I__653 (
            .O(N__4781),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_14 ));
    InMux I__652 (
            .O(N__4776),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_13 ));
    InMux I__651 (
            .O(N__4773),
            .I(N__4769));
    InMux I__650 (
            .O(N__4772),
            .I(N__4766));
    LocalMux I__649 (
            .O(N__4769),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_15 ));
    LocalMux I__648 (
            .O(N__4766),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_15 ));
    InMux I__647 (
            .O(N__4761),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_14 ));
    InMux I__646 (
            .O(N__4758),
            .I(N__4754));
    InMux I__645 (
            .O(N__4757),
            .I(N__4751));
    LocalMux I__644 (
            .O(N__4754),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_16 ));
    LocalMux I__643 (
            .O(N__4751),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_16 ));
    InMux I__642 (
            .O(N__4746),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_15 ));
    InMux I__641 (
            .O(N__4743),
            .I(N__4739));
    InMux I__640 (
            .O(N__4742),
            .I(N__4736));
    LocalMux I__639 (
            .O(N__4739),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_17 ));
    LocalMux I__638 (
            .O(N__4736),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_17 ));
    InMux I__637 (
            .O(N__4731),
            .I(bfn_5_6_0_));
    CascadeMux I__636 (
            .O(N__4728),
            .I(N__4724));
    InMux I__635 (
            .O(N__4727),
            .I(N__4721));
    InMux I__634 (
            .O(N__4724),
            .I(N__4718));
    LocalMux I__633 (
            .O(N__4721),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_18 ));
    LocalMux I__632 (
            .O(N__4718),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_18 ));
    InMux I__631 (
            .O(N__4713),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_17 ));
    InMux I__630 (
            .O(N__4710),
            .I(N__4706));
    InMux I__629 (
            .O(N__4709),
            .I(N__4703));
    LocalMux I__628 (
            .O(N__4706),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_19 ));
    LocalMux I__627 (
            .O(N__4703),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_19 ));
    InMux I__626 (
            .O(N__4698),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_18 ));
    InMux I__625 (
            .O(N__4695),
            .I(N__4691));
    InMux I__624 (
            .O(N__4694),
            .I(N__4688));
    LocalMux I__623 (
            .O(N__4691),
            .I(N__4685));
    LocalMux I__622 (
            .O(N__4688),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_20 ));
    Odrv4 I__621 (
            .O(N__4685),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_20 ));
    InMux I__620 (
            .O(N__4680),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_19 ));
    InMux I__619 (
            .O(N__4677),
            .I(N__4673));
    InMux I__618 (
            .O(N__4676),
            .I(N__4670));
    LocalMux I__617 (
            .O(N__4673),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_21 ));
    LocalMux I__616 (
            .O(N__4670),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_21 ));
    InMux I__615 (
            .O(N__4665),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_20 ));
    CascadeMux I__614 (
            .O(N__4662),
            .I(N__4658));
    InMux I__613 (
            .O(N__4661),
            .I(N__4655));
    InMux I__612 (
            .O(N__4658),
            .I(N__4652));
    LocalMux I__611 (
            .O(N__4655),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_22 ));
    LocalMux I__610 (
            .O(N__4652),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_22 ));
    InMux I__609 (
            .O(N__4647),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_21 ));
    InMux I__608 (
            .O(N__4644),
            .I(N__4640));
    InMux I__607 (
            .O(N__4643),
            .I(N__4637));
    LocalMux I__606 (
            .O(N__4640),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_6 ));
    LocalMux I__605 (
            .O(N__4637),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_6 ));
    InMux I__604 (
            .O(N__4632),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_5 ));
    InMux I__603 (
            .O(N__4629),
            .I(N__4625));
    InMux I__602 (
            .O(N__4628),
            .I(N__4622));
    LocalMux I__601 (
            .O(N__4625),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_7 ));
    LocalMux I__600 (
            .O(N__4622),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_7 ));
    InMux I__599 (
            .O(N__4617),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_6 ));
    CascadeMux I__598 (
            .O(N__4614),
            .I(N__4610));
    InMux I__597 (
            .O(N__4613),
            .I(N__4607));
    InMux I__596 (
            .O(N__4610),
            .I(N__4604));
    LocalMux I__595 (
            .O(N__4607),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_8 ));
    LocalMux I__594 (
            .O(N__4604),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_8 ));
    InMux I__593 (
            .O(N__4599),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_7 ));
    CascadeMux I__592 (
            .O(N__4596),
            .I(N__4592));
    InMux I__591 (
            .O(N__4595),
            .I(N__4589));
    InMux I__590 (
            .O(N__4592),
            .I(N__4586));
    LocalMux I__589 (
            .O(N__4589),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_9 ));
    LocalMux I__588 (
            .O(N__4586),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_9 ));
    InMux I__587 (
            .O(N__4581),
            .I(bfn_5_5_0_));
    InMux I__586 (
            .O(N__4578),
            .I(N__4574));
    InMux I__585 (
            .O(N__4577),
            .I(N__4571));
    LocalMux I__584 (
            .O(N__4574),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_10 ));
    LocalMux I__583 (
            .O(N__4571),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_10 ));
    InMux I__582 (
            .O(N__4566),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_9 ));
    InMux I__581 (
            .O(N__4563),
            .I(N__4559));
    InMux I__580 (
            .O(N__4562),
            .I(N__4556));
    LocalMux I__579 (
            .O(N__4559),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_11 ));
    LocalMux I__578 (
            .O(N__4556),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_11 ));
    InMux I__577 (
            .O(N__4551),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_10 ));
    InMux I__576 (
            .O(N__4548),
            .I(N__4544));
    InMux I__575 (
            .O(N__4547),
            .I(N__4541));
    LocalMux I__574 (
            .O(N__4544),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_12 ));
    LocalMux I__573 (
            .O(N__4541),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_12 ));
    InMux I__572 (
            .O(N__4536),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_11 ));
    InMux I__571 (
            .O(N__4533),
            .I(N__4529));
    InMux I__570 (
            .O(N__4532),
            .I(N__4526));
    LocalMux I__569 (
            .O(N__4529),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_13 ));
    LocalMux I__568 (
            .O(N__4526),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_13 ));
    InMux I__567 (
            .O(N__4521),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_12 ));
    IoInMux I__566 (
            .O(N__4518),
            .I(N__4515));
    LocalMux I__565 (
            .O(N__4515),
            .I(N__4512));
    IoSpan4Mux I__564 (
            .O(N__4512),
            .I(N__4509));
    Odrv4 I__563 (
            .O(N__4509),
            .I(r_Hex_Encoding_i_6));
    IoInMux I__562 (
            .O(N__4506),
            .I(N__4503));
    LocalMux I__561 (
            .O(N__4503),
            .I(r_Hex_Encoding_i_3));
    IoInMux I__560 (
            .O(N__4500),
            .I(N__4497));
    LocalMux I__559 (
            .O(N__4497),
            .I(r_Hex_Encoding_i_0));
    IoInMux I__558 (
            .O(N__4494),
            .I(N__4491));
    LocalMux I__557 (
            .O(N__4491),
            .I(r_Hex_Encoding_i_4));
    InMux I__556 (
            .O(N__4488),
            .I(N__4484));
    InMux I__555 (
            .O(N__4487),
            .I(N__4481));
    LocalMux I__554 (
            .O(N__4484),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_2 ));
    LocalMux I__553 (
            .O(N__4481),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_2 ));
    InMux I__552 (
            .O(N__4476),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_1 ));
    InMux I__551 (
            .O(N__4473),
            .I(N__4469));
    InMux I__550 (
            .O(N__4472),
            .I(N__4466));
    LocalMux I__549 (
            .O(N__4469),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_3 ));
    LocalMux I__548 (
            .O(N__4466),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_3 ));
    InMux I__547 (
            .O(N__4461),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_2 ));
    InMux I__546 (
            .O(N__4458),
            .I(N__4455));
    LocalMux I__545 (
            .O(N__4455),
            .I(N__4451));
    InMux I__544 (
            .O(N__4454),
            .I(N__4448));
    Span4Mux_v I__543 (
            .O(N__4451),
            .I(N__4445));
    LocalMux I__542 (
            .O(N__4448),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_4 ));
    Odrv4 I__541 (
            .O(N__4445),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_4 ));
    InMux I__540 (
            .O(N__4440),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_3 ));
    InMux I__539 (
            .O(N__4437),
            .I(N__4433));
    InMux I__538 (
            .O(N__4436),
            .I(N__4430));
    LocalMux I__537 (
            .O(N__4433),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_5 ));
    LocalMux I__536 (
            .O(N__4430),
            .I(\Game_Inst.Count_Inst.r_CounterZ0Z_5 ));
    InMux I__535 (
            .O(N__4425),
            .I(\Game_Inst.Count_Inst.un3_r_Counter_cry_4 ));
    CascadeMux I__534 (
            .O(N__4422),
            .I(N__4419));
    InMux I__533 (
            .O(N__4419),
            .I(N__4416));
    LocalMux I__532 (
            .O(N__4416),
            .I(\Game_Inst.r_SM_Main_ns_i_m2_ns_1_0 ));
    CascadeMux I__531 (
            .O(N__4413),
            .I(\Game_Inst.N_260_0_cascade_ ));
    CascadeMux I__530 (
            .O(N__4410),
            .I(N__4407));
    InMux I__529 (
            .O(N__4407),
            .I(N__4404));
    LocalMux I__528 (
            .O(N__4404),
            .I(N__4401));
    Odrv4 I__527 (
            .O(N__4401),
            .I(\Game_Inst.N_260_0 ));
    IoInMux I__526 (
            .O(N__4398),
            .I(N__4395));
    LocalMux I__525 (
            .O(N__4395),
            .I(N__4392));
    Odrv12 I__524 (
            .O(N__4392),
            .I(r_Hex_Encoding_i_1));
    IoInMux I__523 (
            .O(N__4389),
            .I(N__4386));
    LocalMux I__522 (
            .O(N__4386),
            .I(N__4383));
    Span4Mux_s1_v I__521 (
            .O(N__4383),
            .I(N__4380));
    Odrv4 I__520 (
            .O(N__4380),
            .I(r_Hex_Encoding_i_5));
    InMux I__519 (
            .O(N__4377),
            .I(N__4374));
    LocalMux I__518 (
            .O(N__4374),
            .I(\Game_Inst.Count_Inst.o_Toggle3_17 ));
    InMux I__517 (
            .O(N__4371),
            .I(N__4365));
    InMux I__516 (
            .O(N__4370),
            .I(N__4365));
    LocalMux I__515 (
            .O(N__4365),
            .I(\Game_Inst.Count_Inst.o_Toggle3_21 ));
    CascadeMux I__514 (
            .O(N__4362),
            .I(\Game_Inst.Count_Inst.o_Toggle3_17_cascade_ ));
    InMux I__513 (
            .O(N__4359),
            .I(N__4353));
    InMux I__512 (
            .O(N__4358),
            .I(N__4353));
    LocalMux I__511 (
            .O(N__4353),
            .I(\Game_Inst.Count_Inst.o_Toggle3_16 ));
    InMux I__510 (
            .O(N__4350),
            .I(N__4347));
    LocalMux I__509 (
            .O(N__4347),
            .I(\Game_Inst.N_249_0 ));
    CascadeMux I__508 (
            .O(N__4344),
            .I(\Game_Inst.Count_Inst.o_Toggle3_cascade_ ));
    CascadeMux I__507 (
            .O(N__4341),
            .I(\Game_Inst.r_SM_Main_ns_i_0_0_cascade_ ));
    CascadeMux I__506 (
            .O(N__4338),
            .I(\Game_Inst.r_SM_Main_ns_i_1_0_cascade_ ));
    CascadeMux I__505 (
            .O(N__4335),
            .I(\Game_Inst.r_SM_Main_ns_i_2_0_cascade_ ));
    InMux I__504 (
            .O(N__4332),
            .I(N__4329));
    LocalMux I__503 (
            .O(N__4329),
            .I(\Game_Inst.N_338 ));
    InMux I__502 (
            .O(N__4326),
            .I(N__4323));
    LocalMux I__501 (
            .O(N__4323),
            .I(\Game_Inst.Count_Inst.o_Toggle3_14 ));
    CascadeMux I__500 (
            .O(N__4320),
            .I(\Game_Inst.Count_Inst.o_Toggle3_13_cascade_ ));
    InMux I__499 (
            .O(N__4317),
            .I(N__4314));
    LocalMux I__498 (
            .O(N__4314),
            .I(\Game_Inst.Count_Inst.o_Toggle3_12 ));
    InMux I__497 (
            .O(N__4311),
            .I(N__4308));
    LocalMux I__496 (
            .O(N__4308),
            .I(\Game_Inst.Count_Inst.o_Toggle3_15 ));
    CascadeMux I__495 (
            .O(N__4305),
            .I(\Game_Inst.N_334_0_cascade_ ));
    CascadeMux I__494 (
            .O(N__4302),
            .I(\Game_Inst.N_249_0_cascade_ ));
    IoInMux I__493 (
            .O(N__4299),
            .I(N__4296));
    LocalMux I__492 (
            .O(N__4296),
            .I(N__4293));
    Span4Mux_s3_h I__491 (
            .O(N__4293),
            .I(N__4290));
    Odrv4 I__490 (
            .O(N__4290),
            .I(\Game_Inst.Count_Inst.r_Counter_RNIGDO97Z0Z_16 ));
    InMux I__489 (
            .O(N__4287),
            .I(bfn_1_13_0_));
    CascadeMux I__488 (
            .O(N__4284),
            .I(N__4281));
    InMux I__487 (
            .O(N__4281),
            .I(N__4276));
    InMux I__486 (
            .O(N__4280),
            .I(N__4272));
    InMux I__485 (
            .O(N__4279),
            .I(N__4269));
    LocalMux I__484 (
            .O(N__4276),
            .I(N__4266));
    InMux I__483 (
            .O(N__4275),
            .I(N__4263));
    LocalMux I__482 (
            .O(N__4272),
            .I(\Debounce_SW1.r_CountZ0Z_0 ));
    LocalMux I__481 (
            .O(N__4269),
            .I(\Debounce_SW1.r_CountZ0Z_0 ));
    Odrv4 I__480 (
            .O(N__4266),
            .I(\Debounce_SW1.r_CountZ0Z_0 ));
    LocalMux I__479 (
            .O(N__4263),
            .I(\Debounce_SW1.r_CountZ0Z_0 ));
    SRMux I__478 (
            .O(N__4254),
            .I(N__4239));
    SRMux I__477 (
            .O(N__4253),
            .I(N__4239));
    SRMux I__476 (
            .O(N__4252),
            .I(N__4239));
    SRMux I__475 (
            .O(N__4251),
            .I(N__4239));
    SRMux I__474 (
            .O(N__4250),
            .I(N__4239));
    GlobalMux I__473 (
            .O(N__4239),
            .I(N__4236));
    gio2CtrlBuf I__472 (
            .O(N__4236),
            .I(\Debounce_SW1.r_Count12_i_g ));
    InMux I__471 (
            .O(N__4233),
            .I(N__4228));
    InMux I__470 (
            .O(N__4232),
            .I(N__4225));
    InMux I__469 (
            .O(N__4231),
            .I(N__4222));
    LocalMux I__468 (
            .O(N__4228),
            .I(N__4219));
    LocalMux I__467 (
            .O(N__4225),
            .I(N__4216));
    LocalMux I__466 (
            .O(N__4222),
            .I(\Debounce_SW1.r_CountZ0Z_17 ));
    Odrv4 I__465 (
            .O(N__4219),
            .I(\Debounce_SW1.r_CountZ0Z_17 ));
    Odrv4 I__464 (
            .O(N__4216),
            .I(\Debounce_SW1.r_CountZ0Z_17 ));
    CascadeMux I__463 (
            .O(N__4209),
            .I(N__4204));
    CascadeMux I__462 (
            .O(N__4208),
            .I(N__4201));
    InMux I__461 (
            .O(N__4207),
            .I(N__4198));
    InMux I__460 (
            .O(N__4204),
            .I(N__4195));
    InMux I__459 (
            .O(N__4201),
            .I(N__4192));
    LocalMux I__458 (
            .O(N__4198),
            .I(\Debounce_SW1.r_CountZ0Z_7 ));
    LocalMux I__457 (
            .O(N__4195),
            .I(\Debounce_SW1.r_CountZ0Z_7 ));
    LocalMux I__456 (
            .O(N__4192),
            .I(\Debounce_SW1.r_CountZ0Z_7 ));
    InMux I__455 (
            .O(N__4185),
            .I(N__4182));
    LocalMux I__454 (
            .O(N__4182),
            .I(\Debounce_SW1.r_Count13_10 ));
    CascadeMux I__453 (
            .O(N__4179),
            .I(\Debounce_SW1.r_Count13_0_a7_4_cascade_ ));
    InMux I__452 (
            .O(N__4176),
            .I(N__4171));
    InMux I__451 (
            .O(N__4175),
            .I(N__4168));
    InMux I__450 (
            .O(N__4174),
            .I(N__4165));
    LocalMux I__449 (
            .O(N__4171),
            .I(\Debounce_SW1.r_CountZ0Z_5 ));
    LocalMux I__448 (
            .O(N__4168),
            .I(\Debounce_SW1.r_CountZ0Z_5 ));
    LocalMux I__447 (
            .O(N__4165),
            .I(\Debounce_SW1.r_CountZ0Z_5 ));
    InMux I__446 (
            .O(N__4158),
            .I(N__4154));
    InMux I__445 (
            .O(N__4157),
            .I(N__4151));
    LocalMux I__444 (
            .O(N__4154),
            .I(N__4146));
    LocalMux I__443 (
            .O(N__4151),
            .I(N__4146));
    Sp12to4 I__442 (
            .O(N__4146),
            .I(N__4143));
    Span12Mux_v I__441 (
            .O(N__4143),
            .I(N__4140));
    Odrv12 I__440 (
            .O(N__4140),
            .I(i_Switch_1_c));
    InMux I__439 (
            .O(N__4137),
            .I(N__4134));
    LocalMux I__438 (
            .O(N__4134),
            .I(\Debounce_SW1.r_Count13_0_a7_7 ));
    CascadeMux I__437 (
            .O(N__4131),
            .I(\Debounce_SW1.r_Count13_0_a7_8_cascade_ ));
    InMux I__436 (
            .O(N__4128),
            .I(N__4123));
    CascadeMux I__435 (
            .O(N__4127),
            .I(N__4120));
    InMux I__434 (
            .O(N__4126),
            .I(N__4117));
    LocalMux I__433 (
            .O(N__4123),
            .I(N__4114));
    InMux I__432 (
            .O(N__4120),
            .I(N__4111));
    LocalMux I__431 (
            .O(N__4117),
            .I(\Debounce_SW1.r_CountZ0Z_16 ));
    Odrv4 I__430 (
            .O(N__4114),
            .I(\Debounce_SW1.r_CountZ0Z_16 ));
    LocalMux I__429 (
            .O(N__4111),
            .I(\Debounce_SW1.r_CountZ0Z_16 ));
    InMux I__428 (
            .O(N__4104),
            .I(N__4100));
    InMux I__427 (
            .O(N__4103),
            .I(N__4096));
    LocalMux I__426 (
            .O(N__4100),
            .I(N__4093));
    InMux I__425 (
            .O(N__4099),
            .I(N__4090));
    LocalMux I__424 (
            .O(N__4096),
            .I(\Debounce_SW1.r_CountZ0Z_12 ));
    Odrv4 I__423 (
            .O(N__4093),
            .I(\Debounce_SW1.r_CountZ0Z_12 ));
    LocalMux I__422 (
            .O(N__4090),
            .I(\Debounce_SW1.r_CountZ0Z_12 ));
    InMux I__421 (
            .O(N__4083),
            .I(N__4080));
    LocalMux I__420 (
            .O(N__4080),
            .I(\Debounce_SW1.un1_r_Count_8lto17_i_2 ));
    InMux I__419 (
            .O(N__4077),
            .I(N__4072));
    InMux I__418 (
            .O(N__4076),
            .I(N__4067));
    InMux I__417 (
            .O(N__4075),
            .I(N__4067));
    LocalMux I__416 (
            .O(N__4072),
            .I(\Debounce_SW1.r_CountZ0Z_15 ));
    LocalMux I__415 (
            .O(N__4067),
            .I(\Debounce_SW1.r_CountZ0Z_15 ));
    InMux I__414 (
            .O(N__4062),
            .I(N__4057));
    InMux I__413 (
            .O(N__4061),
            .I(N__4054));
    InMux I__412 (
            .O(N__4060),
            .I(N__4051));
    LocalMux I__411 (
            .O(N__4057),
            .I(N__4048));
    LocalMux I__410 (
            .O(N__4054),
            .I(\Debounce_SW1.r_CountZ0Z_14 ));
    LocalMux I__409 (
            .O(N__4051),
            .I(\Debounce_SW1.r_CountZ0Z_14 ));
    Odrv4 I__408 (
            .O(N__4048),
            .I(\Debounce_SW1.r_CountZ0Z_14 ));
    InMux I__407 (
            .O(N__4041),
            .I(N__4038));
    LocalMux I__406 (
            .O(N__4038),
            .I(\Debounce_SW1.r_Count13_0_a7_0 ));
    InMux I__405 (
            .O(N__4035),
            .I(N__4031));
    InMux I__404 (
            .O(N__4034),
            .I(N__4028));
    LocalMux I__403 (
            .O(N__4031),
            .I(\Debounce_SW1.r_CountZ0Z_10 ));
    LocalMux I__402 (
            .O(N__4028),
            .I(\Debounce_SW1.r_CountZ0Z_10 ));
    InMux I__401 (
            .O(N__4023),
            .I(N__4019));
    InMux I__400 (
            .O(N__4022),
            .I(N__4016));
    LocalMux I__399 (
            .O(N__4019),
            .I(\Debounce_SW1.r_CountZ0Z_9 ));
    LocalMux I__398 (
            .O(N__4016),
            .I(\Debounce_SW1.r_CountZ0Z_9 ));
    InMux I__397 (
            .O(N__4011),
            .I(N__4006));
    InMux I__396 (
            .O(N__4010),
            .I(N__4001));
    InMux I__395 (
            .O(N__4009),
            .I(N__4001));
    LocalMux I__394 (
            .O(N__4006),
            .I(\Debounce_SW1.r_CountZ0Z_13 ));
    LocalMux I__393 (
            .O(N__4001),
            .I(\Debounce_SW1.r_CountZ0Z_13 ));
    InMux I__392 (
            .O(N__3996),
            .I(N__3990));
    InMux I__391 (
            .O(N__3995),
            .I(N__3990));
    LocalMux I__390 (
            .O(N__3990),
            .I(\Debounce_SW1.N_28_2 ));
    InMux I__389 (
            .O(N__3987),
            .I(N__3983));
    InMux I__388 (
            .O(N__3986),
            .I(N__3980));
    LocalMux I__387 (
            .O(N__3983),
            .I(\Debounce_SW1.r_CountZ0Z_8 ));
    LocalMux I__386 (
            .O(N__3980),
            .I(\Debounce_SW1.r_CountZ0Z_8 ));
    InMux I__385 (
            .O(N__3975),
            .I(\Debounce_SW1.r_Count_1_cry_7 ));
    InMux I__384 (
            .O(N__3972),
            .I(bfn_1_12_0_));
    InMux I__383 (
            .O(N__3969),
            .I(\Debounce_SW1.r_Count_1_cry_9 ));
    InMux I__382 (
            .O(N__3966),
            .I(N__3962));
    InMux I__381 (
            .O(N__3965),
            .I(N__3959));
    LocalMux I__380 (
            .O(N__3962),
            .I(N__3956));
    LocalMux I__379 (
            .O(N__3959),
            .I(\Debounce_SW1.r_CountZ0Z_11 ));
    Odrv4 I__378 (
            .O(N__3956),
            .I(\Debounce_SW1.r_CountZ0Z_11 ));
    InMux I__377 (
            .O(N__3951),
            .I(\Debounce_SW1.r_Count_1_cry_10 ));
    InMux I__376 (
            .O(N__3948),
            .I(\Debounce_SW1.r_Count_1_cry_11 ));
    InMux I__375 (
            .O(N__3945),
            .I(\Debounce_SW1.r_Count_1_cry_12 ));
    InMux I__374 (
            .O(N__3942),
            .I(\Debounce_SW1.r_Count_1_cry_13 ));
    InMux I__373 (
            .O(N__3939),
            .I(\Debounce_SW1.r_Count_1_cry_14 ));
    InMux I__372 (
            .O(N__3936),
            .I(\Debounce_SW1.r_Count_1_cry_15 ));
    CascadeMux I__371 (
            .O(N__3933),
            .I(\Debounce_SW1.r_Count13_10_cascade_ ));
    InMux I__370 (
            .O(N__3930),
            .I(N__3927));
    LocalMux I__369 (
            .O(N__3927),
            .I(\Debounce_SW1.N_30 ));
    InMux I__368 (
            .O(N__3924),
            .I(N__3919));
    InMux I__367 (
            .O(N__3923),
            .I(N__3916));
    InMux I__366 (
            .O(N__3922),
            .I(N__3913));
    LocalMux I__365 (
            .O(N__3919),
            .I(N__3910));
    LocalMux I__364 (
            .O(N__3916),
            .I(N__3907));
    LocalMux I__363 (
            .O(N__3913),
            .I(\Debounce_SW1.r_CountZ0Z_1 ));
    Odrv12 I__362 (
            .O(N__3910),
            .I(\Debounce_SW1.r_CountZ0Z_1 ));
    Odrv4 I__361 (
            .O(N__3907),
            .I(\Debounce_SW1.r_CountZ0Z_1 ));
    InMux I__360 (
            .O(N__3900),
            .I(N__3896));
    InMux I__359 (
            .O(N__3899),
            .I(N__3893));
    LocalMux I__358 (
            .O(N__3896),
            .I(\Debounce_SW1.r_CountZ0Z_2 ));
    LocalMux I__357 (
            .O(N__3893),
            .I(\Debounce_SW1.r_CountZ0Z_2 ));
    InMux I__356 (
            .O(N__3888),
            .I(\Debounce_SW1.r_Count_1_cry_1 ));
    CascadeMux I__355 (
            .O(N__3885),
            .I(N__3881));
    InMux I__354 (
            .O(N__3884),
            .I(N__3878));
    InMux I__353 (
            .O(N__3881),
            .I(N__3875));
    LocalMux I__352 (
            .O(N__3878),
            .I(\Debounce_SW1.r_CountZ0Z_3 ));
    LocalMux I__351 (
            .O(N__3875),
            .I(\Debounce_SW1.r_CountZ0Z_3 ));
    InMux I__350 (
            .O(N__3870),
            .I(\Debounce_SW1.r_Count_1_cry_2 ));
    InMux I__349 (
            .O(N__3867),
            .I(N__3862));
    InMux I__348 (
            .O(N__3866),
            .I(N__3857));
    InMux I__347 (
            .O(N__3865),
            .I(N__3857));
    LocalMux I__346 (
            .O(N__3862),
            .I(\Debounce_SW1.r_CountZ0Z_4 ));
    LocalMux I__345 (
            .O(N__3857),
            .I(\Debounce_SW1.r_CountZ0Z_4 ));
    InMux I__344 (
            .O(N__3852),
            .I(\Debounce_SW1.r_Count_1_cry_3 ));
    InMux I__343 (
            .O(N__3849),
            .I(\Debounce_SW1.r_Count_1_cry_4 ));
    InMux I__342 (
            .O(N__3846),
            .I(N__3841));
    InMux I__341 (
            .O(N__3845),
            .I(N__3836));
    InMux I__340 (
            .O(N__3844),
            .I(N__3836));
    LocalMux I__339 (
            .O(N__3841),
            .I(\Debounce_SW1.r_CountZ0Z_6 ));
    LocalMux I__338 (
            .O(N__3836),
            .I(\Debounce_SW1.r_CountZ0Z_6 ));
    InMux I__337 (
            .O(N__3831),
            .I(\Debounce_SW1.r_Count_1_cry_5 ));
    InMux I__336 (
            .O(N__3828),
            .I(\Debounce_SW1.r_Count_1_cry_6 ));
    IoInMux I__335 (
            .O(N__3825),
            .I(N__3822));
    LocalMux I__334 (
            .O(N__3822),
            .I(\Debounce_SW1.r_Count12_i ));
    CascadeMux I__333 (
            .O(N__3819),
            .I(\Debounce_SW1.N_28_1_cascade_ ));
    InMux I__332 (
            .O(N__3816),
            .I(N__3813));
    LocalMux I__331 (
            .O(N__3813),
            .I(\Debounce_SW1.N_28_1 ));
    InMux I__330 (
            .O(N__3810),
            .I(N__3807));
    LocalMux I__329 (
            .O(N__3807),
            .I(\Debounce_SW1.N_28 ));
    InMux I__328 (
            .O(N__3804),
            .I(N__3801));
    LocalMux I__327 (
            .O(N__3801),
            .I(\Debounce_SW1.un1_r_Count_8lto17_i_3 ));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(\Game_Inst.Count_Inst.un3_r_Counter_cry_8 ),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(\Game_Inst.Count_Inst.un3_r_Counter_cry_16 ),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(\Debounce_SW4.r_Count_1_cry_8 ),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\Debounce_SW4.r_Count_1_cry_16 ),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\Debounce_SW3.r_Count_1_cry_8 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\Debounce_SW3.r_Count_1_cry_16 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_6_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_13_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(\Debounce_SW2.r_Count_1_cry_8 ),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(\Debounce_SW2.r_Count_1_cry_16 ),
            .carryinitout(bfn_6_15_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\Debounce_SW1.r_Count_1_cry_8 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(\Debounce_SW1.r_Count_1_cry_16 ),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    ICE_GB \Debounce_SW2.r_State_RNI5LPJ4_0  (
            .USERSIGNALTOGLOBALBUFFER(N__6738),
            .GLOBALBUFFEROUTPUT(\Debounce_SW2.r_Count12_i_g ));
    ICE_GB \Game_Inst.Count_Inst.r_Counter_RNIGDO97_0_16  (
            .USERSIGNALTOGLOBALBUFFER(N__4299),
            .GLOBALBUFFEROUTPUT(\Game_Inst.Count_Inst.N_213_g ));
    ICE_GB \Debounce_SW4.r_State_RNI9SDT2_0  (
            .USERSIGNALTOGLOBALBUFFER(N__6270),
            .GLOBALBUFFEROUTPUT(\Debounce_SW4.r_Count12_i_g ));
    ICE_GB \Debounce_SW3.r_State_RNIQSU81_0  (
            .USERSIGNALTOGLOBALBUFFER(N__8109),
            .GLOBALBUFFEROUTPUT(\Debounce_SW3.r_Count12_i_g ));
    ICE_GB \Debounce_SW1.r_State_RNIGDKU2_0  (
            .USERSIGNALTOGLOBALBUFFER(N__3825),
            .GLOBALBUFFEROUTPUT(\Debounce_SW1.r_Count12_i_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \Debounce_SW1.r_Count_1_LC_1_8_1 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_1_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_1_LC_1_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Debounce_SW1.r_Count_1_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__3922),
            .in2(_gnd_net_),
            .in3(N__4280),
            .lcout(\Debounce_SW1.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8404),
            .ce(),
            .sr(N__4250));
    defparam \Debounce_SW1.r_State_RNIGDKU2_LC_1_9_7 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_RNIGDKU2_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_State_RNIGDKU2_LC_1_9_7 .LUT_INIT=16'b1100001111010111;
    LogicCell40 \Debounce_SW1.r_State_RNIGDKU2_LC_1_9_7  (
            .in0(N__3804),
            .in1(N__4158),
            .in2(N__6103),
            .in3(N__3810),
            .lcout(\Debounce_SW1.r_Count12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIO539_8_LC_1_10_0 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIO539_8_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIO539_8_LC_1_10_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Debounce_SW1.r_Count_RNIO539_8_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__3966),
            .in2(_gnd_net_),
            .in3(N__3986),
            .lcout(\Debounce_SW1.N_28_1 ),
            .ltout(\Debounce_SW1.N_28_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_State_RNO_0_LC_1_10_1 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_RNO_0_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_State_RNO_0_LC_1_10_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Debounce_SW1.r_State_RNO_0_LC_1_10_1  (
            .in0(N__3845),
            .in1(N__3866),
            .in2(N__3819),
            .in3(N__3996),
            .lcout(\Debounce_SW1.r_Count13_0_a7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNI78LD1_7_LC_1_10_2 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNI78LD1_7_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNI78LD1_7_LC_1_10_2 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \Debounce_SW1.r_Count_RNI78LD1_7_LC_1_10_2  (
            .in0(N__3995),
            .in1(N__3816),
            .in2(N__4208),
            .in3(N__3930),
            .lcout(\Debounce_SW1.N_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIR1R61_17_LC_1_10_4 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIR1R61_17_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIR1R61_17_LC_1_10_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \Debounce_SW1.r_Count_RNIR1R61_17_LC_1_10_4  (
            .in0(N__4232),
            .in1(N__4062),
            .in2(_gnd_net_),
            .in3(N__4083),
            .lcout(\Debounce_SW1.un1_r_Count_8lto17_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNI2KFA_1_LC_1_10_6 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNI2KFA_1_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNI2KFA_1_LC_1_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW1.r_Count_RNI2KFA_1_LC_1_10_6  (
            .in0(N__3899),
            .in1(N__4275),
            .in2(N__3885),
            .in3(N__3923),
            .lcout(\Debounce_SW1.r_Count13_10 ),
            .ltout(\Debounce_SW1.r_Count13_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIULBI_4_LC_1_10_7 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIULBI_4_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIULBI_4_LC_1_10_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Debounce_SW1.r_Count_RNIULBI_4_LC_1_10_7  (
            .in0(N__3844),
            .in1(N__4174),
            .in2(N__3933),
            .in3(N__3865),
            .lcout(\Debounce_SW1.N_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_1_cry_1_c_LC_1_11_0 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_1_cry_1_c_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_1_cry_1_c_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_SW1.r_Count_1_cry_1_c_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__3924),
            .in2(N__4284),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\Debounce_SW1.r_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_2_LC_1_11_1 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_2_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_2_LC_1_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_2_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__3900),
            .in2(_gnd_net_),
            .in3(N__3888),
            .lcout(\Debounce_SW1.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_1 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_2 ),
            .clk(N__8406),
            .ce(),
            .sr(N__4252));
    defparam \Debounce_SW1.r_Count_3_LC_1_11_2 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_3_LC_1_11_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_3_LC_1_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_3_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__3884),
            .in2(_gnd_net_),
            .in3(N__3870),
            .lcout(\Debounce_SW1.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_2 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_3 ),
            .clk(N__8406),
            .ce(),
            .sr(N__4252));
    defparam \Debounce_SW1.r_Count_4_LC_1_11_3 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_4_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_4_LC_1_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_4_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__3867),
            .in2(_gnd_net_),
            .in3(N__3852),
            .lcout(\Debounce_SW1.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_3 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_4 ),
            .clk(N__8406),
            .ce(),
            .sr(N__4252));
    defparam \Debounce_SW1.r_Count_5_LC_1_11_4 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_5_LC_1_11_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_5_LC_1_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_5_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__4175),
            .in2(_gnd_net_),
            .in3(N__3849),
            .lcout(\Debounce_SW1.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_4 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_5 ),
            .clk(N__8406),
            .ce(),
            .sr(N__4252));
    defparam \Debounce_SW1.r_Count_6_LC_1_11_5 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_6_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_6_LC_1_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_6_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__3846),
            .in2(_gnd_net_),
            .in3(N__3831),
            .lcout(\Debounce_SW1.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_5 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_6 ),
            .clk(N__8406),
            .ce(),
            .sr(N__4252));
    defparam \Debounce_SW1.r_Count_7_LC_1_11_6 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_7_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_7_LC_1_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_7_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(N__4207),
            .in2(_gnd_net_),
            .in3(N__3828),
            .lcout(\Debounce_SW1.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_6 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_7 ),
            .clk(N__8406),
            .ce(),
            .sr(N__4252));
    defparam \Debounce_SW1.r_Count_8_LC_1_11_7 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_8_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_8_LC_1_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_8_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__3987),
            .in2(_gnd_net_),
            .in3(N__3975),
            .lcout(\Debounce_SW1.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_7 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_8 ),
            .clk(N__8406),
            .ce(),
            .sr(N__4252));
    defparam \Debounce_SW1.r_Count_9_LC_1_12_0 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_9_LC_1_12_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_9_LC_1_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_9_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__4023),
            .in2(_gnd_net_),
            .in3(N__3972),
            .lcout(\Debounce_SW1.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(\Debounce_SW1.r_Count_1_cry_9 ),
            .clk(N__8409),
            .ce(),
            .sr(N__4253));
    defparam \Debounce_SW1.r_Count_10_LC_1_12_1 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_10_LC_1_12_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_10_LC_1_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_10_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__4035),
            .in2(_gnd_net_),
            .in3(N__3969),
            .lcout(\Debounce_SW1.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_9 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_10 ),
            .clk(N__8409),
            .ce(),
            .sr(N__4253));
    defparam \Debounce_SW1.r_Count_11_LC_1_12_2 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_11_LC_1_12_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_11_LC_1_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_11_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__3965),
            .in2(_gnd_net_),
            .in3(N__3951),
            .lcout(\Debounce_SW1.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_10 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_11 ),
            .clk(N__8409),
            .ce(),
            .sr(N__4253));
    defparam \Debounce_SW1.r_Count_12_LC_1_12_3 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_12_LC_1_12_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_12_LC_1_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_12_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__4103),
            .in2(_gnd_net_),
            .in3(N__3948),
            .lcout(\Debounce_SW1.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_11 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_12 ),
            .clk(N__8409),
            .ce(),
            .sr(N__4253));
    defparam \Debounce_SW1.r_Count_13_LC_1_12_4 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_13_LC_1_12_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_13_LC_1_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_13_LC_1_12_4  (
            .in0(_gnd_net_),
            .in1(N__4011),
            .in2(_gnd_net_),
            .in3(N__3945),
            .lcout(\Debounce_SW1.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_12 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_13 ),
            .clk(N__8409),
            .ce(),
            .sr(N__4253));
    defparam \Debounce_SW1.r_Count_14_LC_1_12_5 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_14_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_14_LC_1_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_14_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__4061),
            .in2(_gnd_net_),
            .in3(N__3942),
            .lcout(\Debounce_SW1.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_13 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_14 ),
            .clk(N__8409),
            .ce(),
            .sr(N__4253));
    defparam \Debounce_SW1.r_Count_15_LC_1_12_6 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_15_LC_1_12_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_15_LC_1_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_15_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__4077),
            .in2(_gnd_net_),
            .in3(N__3939),
            .lcout(\Debounce_SW1.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_14 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_15 ),
            .clk(N__8409),
            .ce(),
            .sr(N__4253));
    defparam \Debounce_SW1.r_Count_16_LC_1_12_7 .C_ON=1'b1;
    defparam \Debounce_SW1.r_Count_16_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_16_LC_1_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW1.r_Count_16_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(N__4126),
            .in2(_gnd_net_),
            .in3(N__3936),
            .lcout(\Debounce_SW1.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_SW1.r_Count_1_cry_15 ),
            .carryout(\Debounce_SW1.r_Count_1_cry_16 ),
            .clk(N__8409),
            .ce(),
            .sr(N__4253));
    defparam \Debounce_SW1.r_Count_17_LC_1_13_0 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_17_LC_1_13_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_17_LC_1_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_SW1.r_Count_17_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__4231),
            .in2(_gnd_net_),
            .in3(N__4287),
            .lcout(\Debounce_SW1.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8413),
            .ce(),
            .sr(N__4254));
    defparam \Debounce_SW1.r_Count_0_LC_2_9_1 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_0_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_Count_0_LC_2_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_SW1.r_Count_0_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4279),
            .lcout(\Debounce_SW1.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8405),
            .ce(),
            .sr(N__4251));
    defparam \Debounce_SW1.r_State_RNO_3_LC_2_10_4 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_RNO_3_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_State_RNO_3_LC_2_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW1.r_State_RNO_3_LC_2_10_4  (
            .in0(N__4128),
            .in1(N__4233),
            .in2(N__4209),
            .in3(N__4104),
            .lcout(),
            .ltout(\Debounce_SW1.r_Count13_0_a7_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_State_RNO_1_LC_2_10_5 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_RNO_1_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_State_RNO_1_LC_2_10_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Debounce_SW1.r_State_RNO_1_LC_2_10_5  (
            .in0(N__4185),
            .in1(N__4041),
            .in2(N__4179),
            .in3(N__4176),
            .lcout(),
            .ltout(\Debounce_SW1.r_Count13_0_a7_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_State_LC_2_10_6 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW1.r_State_LC_2_10_6 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Debounce_SW1.r_State_LC_2_10_6  (
            .in0(N__4157),
            .in1(N__4137),
            .in2(N__4131),
            .in3(N__6086),
            .lcout(w_Switch_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8407),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIGKSP_12_LC_2_11_1 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIGKSP_12_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIGKSP_12_LC_2_11_1 .LUT_INIT=16'b0101111101111111;
    LogicCell40 \Debounce_SW1.r_Count_RNIGKSP_12_LC_2_11_1  (
            .in0(N__4075),
            .in1(N__4009),
            .in2(N__4127),
            .in3(N__4099),
            .lcout(\Debounce_SW1.un1_r_Count_8lto17_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_State_RNO_2_LC_2_11_3 .C_ON=1'b0;
    defparam \Debounce_SW1.r_State_RNO_2_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_State_RNO_2_LC_2_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Debounce_SW1.r_State_RNO_2_LC_2_11_3  (
            .in0(N__4076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4060),
            .lcout(\Debounce_SW1.r_Count13_0_a7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW1.r_Count_RNIR9IF_9_LC_2_11_7 .C_ON=1'b0;
    defparam \Debounce_SW1.r_Count_RNIR9IF_9_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW1.r_Count_RNIR9IF_9_LC_2_11_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Debounce_SW1.r_Count_RNIR9IF_9_LC_2_11_7  (
            .in0(N__4034),
            .in1(N__4022),
            .in2(_gnd_net_),
            .in3(N__4010),
            .lcout(\Debounce_SW1.N_28_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNIN50N1_1_LC_4_4_5 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIN50N1_1_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIN50N1_1_LC_4_4_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNIN50N1_1_LC_4_4_5  (
            .in0(N__4472),
            .in1(N__5148),
            .in2(N__4596),
            .in3(N__4487),
            .lcout(\Game_Inst.Count_Inst.o_Toggle3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNI2H0N1_5_LC_4_4_6 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI2H0N1_5_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI2H0N1_5_LC_4_4_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNI2H0N1_5_LC_4_4_6  (
            .in0(N__4628),
            .in1(N__4643),
            .in2(N__4614),
            .in3(N__4436),
            .lcout(\Game_Inst.Count_Inst.o_Toggle3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNIQ8NM_23_LC_4_5_2 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIQ8NM_23_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIQ8NM_23_LC_4_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNIQ8NM_23_LC_4_5_2  (
            .in0(N__4676),
            .in1(N__4772),
            .in2(N__4833),
            .in3(N__4532),
            .lcout(),
            .ltout(\Game_Inst.Count_Inst.o_Toggle3_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNI6VCR4_10_LC_4_5_3 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI6VCR4_10_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNI6VCR4_10_LC_4_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNI6VCR4_10_LC_4_5_3  (
            .in0(N__4311),
            .in1(N__4326),
            .in2(N__4320),
            .in3(N__4317),
            .lcout(\Game_Inst.Count_Inst.o_Toggle3_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNIJVKM_10_LC_4_5_7 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIJVKM_10_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIJVKM_10_LC_4_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNIJVKM_10_LC_4_5_7  (
            .in0(N__4547),
            .in1(N__4562),
            .in2(N__4791),
            .in3(N__4577),
            .lcout(\Game_Inst.Count_Inst.o_Toggle3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI5RM6_1_LC_4_6_0 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI5RM6_1_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI5RM6_1_LC_4_6_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNI5RM6_1_LC_4_6_0  (
            .in0(N__5661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5749),
            .lcout(\Game_Inst.N_334_0 ),
            .ltout(\Game_Inst.N_334_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIE5PG_2_LC_4_6_1 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIE5PG_2_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIE5PG_2_LC_4_6_1 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \Game_Inst.r_SM_Main_RNIE5PG_2_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__5834),
            .in2(N__4305),
            .in3(N__5473),
            .lcout(\Game_Inst.N_249_0 ),
            .ltout(\Game_Inst.N_249_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNIGDO97_16_LC_4_6_2 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIGDO97_16_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIGDO97_16_LC_4_6_2 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNIGDO97_16_LC_4_6_2  (
            .in0(N__4358),
            .in1(N__4377),
            .in2(N__4302),
            .in3(N__4370),
            .lcout(\Game_Inst.Count_Inst.r_Counter_RNIGDO97Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNIANLM_16_LC_4_6_3 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIANLM_16_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIANLM_16_LC_4_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNIANLM_16_LC_4_6_3  (
            .in0(N__4757),
            .in1(N__4709),
            .in2(N__4728),
            .in3(N__4742),
            .lcout(\Game_Inst.Count_Inst.o_Toggle3_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_RNIIHS61_20_LC_4_6_4 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIIHS61_20_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.r_Counter_RNIIHS61_20_LC_4_6_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_RNIIHS61_20_LC_4_6_4  (
            .in0(N__4695),
            .in1(N__4458),
            .in2(N__4662),
            .in3(N__5169),
            .lcout(\Game_Inst.Count_Inst.o_Toggle3_17 ),
            .ltout(\Game_Inst.Count_Inst.o_Toggle3_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.o_Toggle_RNO_0_LC_4_6_5 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.o_Toggle_RNO_0_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.o_Toggle_RNO_0_LC_4_6_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Game_Inst.Count_Inst.o_Toggle_RNO_0_LC_4_6_5  (
            .in0(N__4371),
            .in1(_gnd_net_),
            .in2(N__4362),
            .in3(N__4359),
            .lcout(),
            .ltout(\Game_Inst.Count_Inst.o_Toggle3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.o_Toggle_LC_4_6_6 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.o_Toggle_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.o_Toggle_LC_4_6_6 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \Game_Inst.Count_Inst.o_Toggle_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(N__4350),
            .in2(N__4344),
            .in3(N__4926),
            .lcout(\Game_Inst.w_Toggle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8415),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_4_0_LC_4_7_0 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_4_0_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_4_0_LC_4_7_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_4_0_LC_4_7_0  (
            .in0(N__5747),
            .in1(N__7581),
            .in2(N__5884),
            .in3(N__6113),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_3_0_LC_4_7_1 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_3_0_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_3_0_LC_4_7_1 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_3_0_LC_4_7_1  (
            .in0(N__4885),
            .in1(N__5748),
            .in2(N__4341),
            .in3(N__5655),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_1_0_LC_4_7_2 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_1_0_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_1_0_LC_4_7_2 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_1_0_LC_4_7_2  (
            .in0(N__5657),
            .in1(N__4854),
            .in2(N__4338),
            .in3(N__5872),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_0_LC_4_7_3 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_0_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_SM_Main_0_LC_4_7_3 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Game_Inst.r_SM_Main_0_LC_4_7_3  (
            .in0(N__4332),
            .in1(N__4817),
            .in2(N__4335),
            .in3(N__4866),
            .lcout(\Game_Inst.r_SM_MainZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8410),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI7TM6_1_LC_4_7_4 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI7TM6_1_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI7TM6_1_LC_4_7_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Game_Inst.r_SM_Main_RNI7TM6_1_LC_4_7_4  (
            .in0(N__5746),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5871),
            .lcout(\Game_Inst.r_SM_Main_ns_i_a4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_0_0_LC_4_7_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_0_0_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_0_0_LC_4_7_5 .LUT_INIT=16'b0010001000001111;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_0_0_LC_4_7_5  (
            .in0(N__4902),
            .in1(N__4925),
            .in2(N__4422),
            .in3(N__5656),
            .lcout(\Game_Inst.N_338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI5RM6_0_1_LC_4_7_7 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI5RM6_0_1_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI5RM6_0_1_LC_4_7_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Game_Inst.r_SM_Main_RNI5RM6_0_1_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(N__5745),
            .in2(_gnd_net_),
            .in3(N__5654),
            .lcout(\Game_Inst.N_310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_2_0_LC_4_8_1 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_2_0_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_2_0_LC_4_8_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_2_0_LC_4_8_1  (
            .in0(N__4976),
            .in1(N__7583),
            .in2(_gnd_net_),
            .in3(N__6112),
            .lcout(\Game_Inst.r_SM_Main_ns_i_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_LC_4_9_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_LC_4_9_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Button_DV_LC_4_9_1 .LUT_INIT=16'b1011101111111011;
    LogicCell40 \Game_Inst.r_Button_DV_LC_4_9_1  (
            .in0(N__6513),
            .in1(N__7359),
            .in2(N__6133),
            .in3(N__6108),
            .lcout(\Game_Inst.r_Button_DVZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8411),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_RNI2T5J1_3_LC_4_9_3 .C_ON=1'b0;
    defparam \Game_Inst.o_Score_RNI2T5J1_3_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.o_Score_RNI2T5J1_3_LC_4_9_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Game_Inst.o_Score_RNI2T5J1_3_LC_4_9_3  (
            .in0(N__5425),
            .in1(N__5350),
            .in2(N__5287),
            .in3(N__5221),
            .lcout(\Game_Inst.N_333_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI6HDK_1_LC_4_10_0 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI6HDK_1_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI6HDK_1_LC_4_10_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Game_Inst.r_SM_Main_RNI6HDK_1_LC_4_10_0  (
            .in0(N__5767),
            .in1(N__5886),
            .in2(_gnd_net_),
            .in3(N__6174),
            .lcout(\Game_Inst.N_260_0 ),
            .ltout(\Game_Inst.N_260_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_0_LC_4_10_1 .C_ON=1'b0;
    defparam \Game_Inst.o_Score_0_LC_4_10_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.o_Score_0_LC_4_10_1 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \Game_Inst.o_Score_0_LC_4_10_1  (
            .in0(N__4950),
            .in1(N__5509),
            .in2(N__4413),
            .in3(N__5546),
            .lcout(w_Score_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8414),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_1_LC_4_10_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_1_LC_4_10_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Switch_1_LC_4_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Switch_1_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6090),
            .lcout(\Game_Inst.r_SwitchZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8414),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_2_LC_4_10_7 .C_ON=1'b0;
    defparam \Game_Inst.o_Score_2_LC_4_10_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.o_Score_2_LC_4_10_7 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \Game_Inst.o_Score_2_LC_4_10_7  (
            .in0(N__5510),
            .in1(N__5547),
            .in2(N__4410),
            .in3(N__4941),
            .lcout(w_Score_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8414),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_1_LC_4_12_3 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_1_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_1_LC_4_12_3 .LUT_INIT=16'b0100101100000010;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_1_LC_4_12_3  (
            .in0(N__5439),
            .in1(N__5379),
            .in2(N__5319),
            .in3(N__5241),
            .lcout(r_Hex_Encoding_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8421),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_5_LC_4_15_6 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_5_LC_4_15_6 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_5_LC_4_15_6 .LUT_INIT=16'b1010010011001000;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_5_LC_4_15_6  (
            .in0(N__5453),
            .in1(N__5391),
            .in2(N__5321),
            .in3(N__5242),
            .lcout(r_Hex_Encoding_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8435),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_6_LC_4_16_1 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_6_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_6_LC_4_16_1 .LUT_INIT=16'b0100100100010000;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_6_LC_4_16_1  (
            .in0(N__5457),
            .in1(N__5318),
            .in2(N__5394),
            .in3(N__5246),
            .lcout(r_Hex_Encoding_i_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8442),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_3_LC_4_16_4 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_3_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_3_LC_4_16_4 .LUT_INIT=16'b1000100101000010;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_3_LC_4_16_4  (
            .in0(N__5244),
            .in1(N__5455),
            .in2(N__5322),
            .in3(N__5389),
            .lcout(r_Hex_Encoding_i_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8442),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_0_LC_4_16_5 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_0_LC_4_16_5 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_0_LC_4_16_5 .LUT_INIT=16'b0010000101000001;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_0_LC_4_16_5  (
            .in0(N__5454),
            .in1(N__5316),
            .in2(N__5392),
            .in3(N__5243),
            .lcout(r_Hex_Encoding_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8442),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_4_LC_4_16_7 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_4_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_4_LC_4_16_7 .LUT_INIT=16'b1000000011000010;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_4_LC_4_16_7  (
            .in0(N__5456),
            .in1(N__5317),
            .in2(N__5393),
            .in3(N__5245),
            .lcout(r_Hex_Encoding_i_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8442),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.un3_r_Counter_cry_1_c_LC_5_4_0 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.un3_r_Counter_cry_1_c_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.Count_Inst.un3_r_Counter_cry_1_c_LC_5_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Game_Inst.Count_Inst.un3_r_Counter_cry_1_c_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(N__5146),
            .in2(N__5181),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_2_LC_5_4_1 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_2_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_2_LC_5_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_2_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__4488),
            .in2(_gnd_net_),
            .in3(N__4476),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_2 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_1 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_2 ),
            .clk(N__8426),
            .ce(),
            .sr(N__5126));
    defparam \Game_Inst.Count_Inst.r_Counter_3_LC_5_4_2 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_3_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_3_LC_5_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_3_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__4473),
            .in2(_gnd_net_),
            .in3(N__4461),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_3 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_2 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_3 ),
            .clk(N__8426),
            .ce(),
            .sr(N__5126));
    defparam \Game_Inst.Count_Inst.r_Counter_4_LC_5_4_3 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_4_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_4_LC_5_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_4_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(N__4454),
            .in2(_gnd_net_),
            .in3(N__4440),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_4 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_3 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_4 ),
            .clk(N__8426),
            .ce(),
            .sr(N__5126));
    defparam \Game_Inst.Count_Inst.r_Counter_5_LC_5_4_4 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_5_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_5_LC_5_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_5_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(N__4437),
            .in2(_gnd_net_),
            .in3(N__4425),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_5 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_4 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_5 ),
            .clk(N__8426),
            .ce(),
            .sr(N__5126));
    defparam \Game_Inst.Count_Inst.r_Counter_6_LC_5_4_5 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_6_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_6_LC_5_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_6_LC_5_4_5  (
            .in0(_gnd_net_),
            .in1(N__4644),
            .in2(_gnd_net_),
            .in3(N__4632),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_6 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_5 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_6 ),
            .clk(N__8426),
            .ce(),
            .sr(N__5126));
    defparam \Game_Inst.Count_Inst.r_Counter_7_LC_5_4_6 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_7_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_7_LC_5_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_7_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__4629),
            .in2(_gnd_net_),
            .in3(N__4617),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_7 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_6 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_7 ),
            .clk(N__8426),
            .ce(),
            .sr(N__5126));
    defparam \Game_Inst.Count_Inst.r_Counter_8_LC_5_4_7 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_8_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_8_LC_5_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_8_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(N__4613),
            .in2(_gnd_net_),
            .in3(N__4599),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_8 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_7 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_8 ),
            .clk(N__8426),
            .ce(),
            .sr(N__5126));
    defparam \Game_Inst.Count_Inst.r_Counter_9_LC_5_5_0 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_9_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_9_LC_5_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_9_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(N__4595),
            .in2(_gnd_net_),
            .in3(N__4581),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_5_0_),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_9 ),
            .clk(N__8422),
            .ce(),
            .sr(N__5125));
    defparam \Game_Inst.Count_Inst.r_Counter_10_LC_5_5_1 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_10_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_10_LC_5_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_10_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__4578),
            .in2(_gnd_net_),
            .in3(N__4566),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_10 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_9 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_10 ),
            .clk(N__8422),
            .ce(),
            .sr(N__5125));
    defparam \Game_Inst.Count_Inst.r_Counter_11_LC_5_5_2 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_11_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_11_LC_5_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_11_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__4563),
            .in2(_gnd_net_),
            .in3(N__4551),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_11 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_10 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_11 ),
            .clk(N__8422),
            .ce(),
            .sr(N__5125));
    defparam \Game_Inst.Count_Inst.r_Counter_12_LC_5_5_3 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_12_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_12_LC_5_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_12_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__4548),
            .in2(_gnd_net_),
            .in3(N__4536),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_12 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_11 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_12 ),
            .clk(N__8422),
            .ce(),
            .sr(N__5125));
    defparam \Game_Inst.Count_Inst.r_Counter_13_LC_5_5_4 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_13_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_13_LC_5_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_13_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__4533),
            .in2(_gnd_net_),
            .in3(N__4521),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_13 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_12 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_13 ),
            .clk(N__8422),
            .ce(),
            .sr(N__5125));
    defparam \Game_Inst.Count_Inst.r_Counter_14_LC_5_5_5 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_14_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_14_LC_5_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_14_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(N__4790),
            .in2(_gnd_net_),
            .in3(N__4776),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_14 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_13 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_14 ),
            .clk(N__8422),
            .ce(),
            .sr(N__5125));
    defparam \Game_Inst.Count_Inst.r_Counter_15_LC_5_5_6 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_15_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_15_LC_5_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_15_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(N__4773),
            .in2(_gnd_net_),
            .in3(N__4761),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_15 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_14 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_15 ),
            .clk(N__8422),
            .ce(),
            .sr(N__5125));
    defparam \Game_Inst.Count_Inst.r_Counter_16_LC_5_5_7 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_16_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_16_LC_5_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_16_LC_5_5_7  (
            .in0(_gnd_net_),
            .in1(N__4758),
            .in2(_gnd_net_),
            .in3(N__4746),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_16 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_15 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_16 ),
            .clk(N__8422),
            .ce(),
            .sr(N__5125));
    defparam \Game_Inst.Count_Inst.r_Counter_17_LC_5_6_0 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_17_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_17_LC_5_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_17_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__4743),
            .in2(_gnd_net_),
            .in3(N__4731),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_17 ),
            .clk(N__8419),
            .ce(),
            .sr(N__5124));
    defparam \Game_Inst.Count_Inst.r_Counter_18_LC_5_6_1 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_18_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_18_LC_5_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_18_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__4727),
            .in2(_gnd_net_),
            .in3(N__4713),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_18 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_17 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_18 ),
            .clk(N__8419),
            .ce(),
            .sr(N__5124));
    defparam \Game_Inst.Count_Inst.r_Counter_19_LC_5_6_2 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_19_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_19_LC_5_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_19_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__4710),
            .in2(_gnd_net_),
            .in3(N__4698),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_19 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_18 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_19 ),
            .clk(N__8419),
            .ce(),
            .sr(N__5124));
    defparam \Game_Inst.Count_Inst.r_Counter_20_LC_5_6_3 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_20_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_20_LC_5_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_20_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__4694),
            .in2(_gnd_net_),
            .in3(N__4680),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_20 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_19 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_20 ),
            .clk(N__8419),
            .ce(),
            .sr(N__5124));
    defparam \Game_Inst.Count_Inst.r_Counter_21_LC_5_6_4 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_21_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_21_LC_5_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_21_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(N__4677),
            .in2(_gnd_net_),
            .in3(N__4665),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_21 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_20 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_21 ),
            .clk(N__8419),
            .ce(),
            .sr(N__5124));
    defparam \Game_Inst.Count_Inst.r_Counter_22_LC_5_6_5 .C_ON=1'b1;
    defparam \Game_Inst.Count_Inst.r_Counter_22_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_22_LC_5_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_22_LC_5_6_5  (
            .in0(_gnd_net_),
            .in1(N__4661),
            .in2(_gnd_net_),
            .in3(N__4647),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_22 ),
            .ltout(),
            .carryin(\Game_Inst.Count_Inst.un3_r_Counter_cry_21 ),
            .carryout(\Game_Inst.Count_Inst.un3_r_Counter_cry_22 ),
            .clk(N__8419),
            .ce(),
            .sr(N__5124));
    defparam \Game_Inst.Count_Inst.r_Counter_23_LC_5_6_6 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_23_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_23_LC_5_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_23_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(N__4832),
            .in2(_gnd_net_),
            .in3(N__4836),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8419),
            .ce(),
            .sr(N__5124));
    defparam \Game_Inst.Count_Inst.r_Counter_0_LC_5_6_7 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_0_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_0_LC_5_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_0_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5173),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8419),
            .ce(),
            .sr(N__5124));
    defparam \Game_Inst.r_Toggle_LC_5_7_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Toggle_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Toggle_LC_5_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Toggle_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4924),
            .lcout(\Game_Inst.r_ToggleZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8416),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_2_LC_5_7_1 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_2_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_SM_Main_2_LC_5_7_1 .LUT_INIT=16'b1100110001001100;
    LogicCell40 \Game_Inst.r_SM_Main_2_LC_5_7_1  (
            .in0(N__5922),
            .in1(N__5019),
            .in2(N__5066),
            .in3(N__5010),
            .lcout(\Game_Inst.r_SM_MainZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8416),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_1_1_LC_5_7_2 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_1_1_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_1_1_LC_5_7_2 .LUT_INIT=16'b0010001100001111;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_1_1_LC_5_7_2  (
            .in0(N__4887),
            .in1(N__5876),
            .in2(N__4818),
            .in3(N__5659),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_0_1_LC_5_7_3 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_0_1_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_0_1_LC_5_7_3 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_0_1_LC_5_7_3  (
            .in0(N__4797),
            .in1(N__5031),
            .in2(N__4803),
            .in3(N__5008),
            .lcout(),
            .ltout(\Game_Inst.r_SM_Main_ns_i_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_1_LC_5_7_4 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_1_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_SM_Main_1_LC_5_7_4 .LUT_INIT=16'b0100000011110000;
    LogicCell40 \Game_Inst.r_SM_Main_1_LC_5_7_4  (
            .in0(N__5009),
            .in1(N__5921),
            .in2(N__4800),
            .in3(N__5045),
            .lcout(\Game_Inst.r_SM_MainZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8416),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_2_1_LC_5_7_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_2_1_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_2_1_LC_5_7_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_2_1_LC_5_7_5  (
            .in0(N__5660),
            .in1(_gnd_net_),
            .in2(N__5885),
            .in3(N__4886),
            .lcout(\Game_Inst.r_SM_Main_ns_i_a4_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Toggle_RNI3C1M_LC_5_7_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Toggle_RNI3C1M_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Toggle_RNI3C1M_LC_5_7_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Game_Inst.r_Toggle_RNI3C1M_LC_5_7_6  (
            .in0(N__4900),
            .in1(N__4922),
            .in2(_gnd_net_),
            .in3(N__5658),
            .lcout(\Game_Inst.N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Toggle_RNI1VLI_LC_5_7_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Toggle_RNI1VLI_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Toggle_RNI1VLI_LC_5_7_7 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \Game_Inst.r_Toggle_RNI1VLI_LC_5_7_7  (
            .in0(N__4923),
            .in1(N__4901),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.r_SM_Main7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_RNIG6DF_LC_5_8_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_RNIG6DF_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_DV_RNIG6DF_LC_5_8_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Game_Inst.r_Button_DV_RNIG6DF_LC_5_8_0  (
            .in0(N__5663),
            .in1(N__5750),
            .in2(_gnd_net_),
            .in3(N__4975),
            .lcout(\Game_Inst.r_SM_Main_0_sqmuxa_2_1 ),
            .ltout(\Game_Inst.r_SM_Main_0_sqmuxa_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_RNI2TG99_LC_5_8_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_RNI2TG99_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_DV_RNI2TG99_LC_5_8_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Game_Inst.r_Button_DV_RNI2TG99_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__5000),
            .in2(N__4869),
            .in3(N__5914),
            .lcout(\Game_Inst.N_345 ),
            .ltout(\Game_Inst.N_345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI5SIOD_1_LC_5_8_2 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI5SIOD_1_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI5SIOD_1_LC_5_8_2 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \Game_Inst.r_SM_Main_RNI5SIOD_1_LC_5_8_2  (
            .in0(N__5504),
            .in1(N__6173),
            .in2(N__4860),
            .in3(N__4986),
            .lcout(\Game_Inst.r_Index_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNO_0_1_LC_5_8_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNO_0_1_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNO_0_1_LC_5_8_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \Game_Inst.r_Index_RNO_0_1_LC_5_8_3  (
            .in0(N__5603),
            .in1(N__6003),
            .in2(_gnd_net_),
            .in3(N__6578),
            .lcout(),
            .ltout(\Game_Inst.SUM_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_1_LC_5_8_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_1_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Index_1_LC_5_8_4 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \Game_Inst.r_Index_1_LC_5_8_4  (
            .in0(N__5975),
            .in1(N__5586),
            .in2(N__4857),
            .in3(N__5703),
            .lcout(\Game_Inst.r_IndexZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8408),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_RNIDO1C_LC_5_8_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_RNIDO1C_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_DV_RNIDO1C_LC_5_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Game_Inst.r_Button_DV_RNIDO1C_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(N__4974),
            .in2(_gnd_net_),
            .in3(N__5662),
            .lcout(\Game_Inst.N_311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_RNI6CJ72_3_LC_5_8_7 .C_ON=1'b0;
    defparam \Game_Inst.o_Score_RNI6CJ72_3_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.o_Score_RNI6CJ72_3_LC_5_8_7 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \Game_Inst.o_Score_RNI6CJ72_3_LC_5_8_7  (
            .in0(N__6172),
            .in1(N__4853),
            .in2(_gnd_net_),
            .in3(N__5474),
            .lcout(\Game_Inst.N_335_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNIU4S41_2_LC_5_9_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNIU4S41_2_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNIU4S41_2_LC_5_9_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Game_Inst.r_Index_RNIU4S41_2_LC_5_9_2  (
            .in0(N__5220),
            .in1(N__5961),
            .in2(N__5372),
            .in3(N__6571),
            .lcout(),
            .ltout(\Game_Inst.r_Index16_NE_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNI7O342_1_LC_5_9_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNI7O342_1_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNI7O342_1_LC_5_9_3 .LUT_INIT=16'b0010000000010000;
    LogicCell40 \Game_Inst.r_Index_RNI7O342_1_LC_5_9_3  (
            .in0(N__5424),
            .in1(N__5288),
            .in2(N__5013),
            .in3(N__6001),
            .lcout(\Game_Inst.N_330_li ),
            .ltout(\Game_Inst.N_330_li_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIH1S03_1_LC_5_9_4 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIH1S03_1_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIH1S03_1_LC_5_9_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNIH1S03_1_LC_5_9_4  (
            .in0(N__5766),
            .in1(N__5869),
            .in2(N__4989),
            .in3(N__5788),
            .lcout(\Game_Inst.r_SM_Main_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_1_LC_5_9_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_1_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_0_1_LC_5_9_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Game_Inst.r_SM_Main_RNI9A2A_0_1_LC_5_9_5  (
            .in0(N__5868),
            .in1(N__5765),
            .in2(_gnd_net_),
            .in3(N__5676),
            .lcout(\Game_Inst.r_SM_Main_98_d ),
            .ltout(\Game_Inst.r_SM_Main_98_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_DV_RNIJ9F01_LC_5_9_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_DV_RNIJ9F01_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_DV_RNIJ9F01_LC_5_9_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Game_Inst.r_Button_DV_RNIJ9F01_LC_5_9_6  (
            .in0(N__4977),
            .in1(N__7584),
            .in2(N__4953),
            .in3(N__6107),
            .lcout(\Game_Inst.o_Score_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_RNO_0_0_LC_5_10_0 .C_ON=1'b1;
    defparam \Game_Inst.o_Score_RNO_0_0_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.o_Score_RNO_0_0_LC_5_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.o_Score_RNO_0_0_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__5222),
            .in2(N__5532),
            .in3(N__5530),
            .lcout(\Game_Inst.o_Score_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\Game_Inst.un1_o_Score_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_RNO_0_1_LC_5_10_1 .C_ON=1'b1;
    defparam \Game_Inst.o_Score_RNO_0_1_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.o_Score_RNO_0_1_LC_5_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.o_Score_RNO_0_1_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__5426),
            .in2(_gnd_net_),
            .in3(N__4944),
            .lcout(\Game_Inst.o_Score_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\Game_Inst.un1_o_Score_cry_0 ),
            .carryout(\Game_Inst.un1_o_Score_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_RNO_0_2_LC_5_10_2 .C_ON=1'b1;
    defparam \Game_Inst.o_Score_RNO_0_2_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.o_Score_RNO_0_2_LC_5_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Game_Inst.o_Score_RNO_0_2_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__5354),
            .in2(_gnd_net_),
            .in3(N__4935),
            .lcout(\Game_Inst.o_Score_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\Game_Inst.un1_o_Score_cry_1 ),
            .carryout(\Game_Inst.un1_o_Score_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_RNO_0_3_LC_5_10_3 .C_ON=1'b0;
    defparam \Game_Inst.o_Score_RNO_0_3_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.o_Score_RNO_0_3_LC_5_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Game_Inst.o_Score_RNO_0_3_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__5286),
            .in2(_gnd_net_),
            .in3(N__4932),
            .lcout(),
            .ltout(\Game_Inst.o_Score_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_3_LC_5_10_4 .C_ON=1'b0;
    defparam \Game_Inst.o_Score_3_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.o_Score_3_LC_5_10_4 .LUT_INIT=16'b0011000100110000;
    LogicCell40 \Game_Inst.o_Score_3_LC_5_10_4  (
            .in0(N__5481),
            .in1(N__5508),
            .in2(N__4929),
            .in3(N__5531),
            .lcout(w_Score_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8418),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI332H_2_LC_5_10_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI332H_2_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI332H_2_LC_5_10_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Game_Inst.r_SM_Main_RNI332H_2_LC_5_10_5  (
            .in0(N__5870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6163),
            .lcout(\Game_Inst.N_287_0 ),
            .ltout(\Game_Inst.N_287_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI5GDK_0_LC_5_10_6 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI5GDK_0_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI5GDK_0_LC_5_10_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNI5GDK_0_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5550),
            .in3(N__5677),
            .lcout(\Game_Inst.N_262_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.o_Score_1_LC_5_10_7 .C_ON=1'b0;
    defparam \Game_Inst.o_Score_1_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.o_Score_1_LC_5_10_7 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \Game_Inst.o_Score_1_LC_5_10_7  (
            .in0(N__5538),
            .in1(N__5529),
            .in2(N__5511),
            .in3(N__5480),
            .lcout(w_Score_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8418),
            .ce(),
            .sr(_gnd_net_));
    defparam \Scoreboard.r_Hex_Encoding_i_2_LC_5_16_6 .C_ON=1'b0;
    defparam \Scoreboard.r_Hex_Encoding_i_2_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \Scoreboard.r_Hex_Encoding_i_2_LC_5_16_6 .LUT_INIT=16'b0001111100000100;
    LogicCell40 \Scoreboard.r_Hex_Encoding_i_2_LC_5_16_6  (
            .in0(N__5452),
            .in1(N__5390),
            .in2(N__5320),
            .in3(N__5250),
            .lcout(r_Hex_Encoding_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8445),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.Count_Inst.r_Counter_1_LC_6_4_0 .C_ON=1'b0;
    defparam \Game_Inst.Count_Inst.r_Counter_1_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.Count_Inst.r_Counter_1_LC_6_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Game_Inst.Count_Inst.r_Counter_1_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__5180),
            .in2(_gnd_net_),
            .in3(N__5147),
            .lcout(\Game_Inst.Count_Inst.r_CounterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8429),
            .ce(),
            .sr(N__5127));
    defparam \Game_Inst.r_SM_Main_RNI9A2A_1_LC_6_7_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_1_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI9A2A_1_LC_6_7_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Game_Inst.r_SM_Main_RNI9A2A_1_LC_6_7_5  (
            .in0(N__5764),
            .in1(N__5866),
            .in2(_gnd_net_),
            .in3(N__5681),
            .lcout(\Game_Inst.r_SM_Main_100_d ),
            .ltout(\Game_Inst.r_SM_Main_100_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI6V986_1_LC_6_7_6 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI6V986_1_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI6V986_1_LC_6_7_6 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \Game_Inst.r_SM_Main_RNI6V986_1_LC_6_7_6  (
            .in0(N__7874),
            .in1(N__6114),
            .in2(N__5085),
            .in3(N__7907),
            .lcout(Game_Inst_o_LED_1_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNO_0_2_LC_6_7_7 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNO_0_2_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNO_0_2_LC_6_7_7 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNO_0_2_LC_6_7_7  (
            .in0(N__5067),
            .in1(N__5865),
            .in2(N__5046),
            .in3(N__5030),
            .lcout(\Game_Inst.r_SM_Main_ns_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNIDV7G1_1_LC_6_8_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNIDV7G1_1_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNIDV7G1_1_LC_6_8_0 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \Game_Inst.r_Index_RNIDV7G1_1_LC_6_8_0  (
            .in0(N__5956),
            .in1(N__5999),
            .in2(N__6309),
            .in3(N__6300),
            .lcout(\Game_Inst.un1_r_Pattern_0__7_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_2__RNIFHRI_0_LC_6_8_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_2__RNIFHRI_0_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_2__RNIFHRI_0_LC_6_8_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Game_Inst.r_Pattern_2__RNIFHRI_0_LC_6_8_1  (
            .in0(N__6562),
            .in1(N__6381),
            .in2(_gnd_net_),
            .in3(N__6375),
            .lcout(\Game_Inst.r_Pattern_2__RNIFHRIZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_0_LC_6_8_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_0_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Index_0_LC_6_8_2 .LUT_INIT=16'b0001010100010000;
    LogicCell40 \Game_Inst.r_Index_0_LC_6_8_2  (
            .in0(N__5585),
            .in1(N__5702),
            .in2(N__6582),
            .in3(N__5604),
            .lcout(\Game_Inst.r_IndexZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8412),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI31SF8_0_LC_6_8_3 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI31SF8_0_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI31SF8_0_LC_6_8_3 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \Game_Inst.r_SM_Main_RNI31SF8_0_LC_6_8_3  (
            .in0(N__5682),
            .in1(N__5562),
            .in2(N__5883),
            .in3(N__5915),
            .lcout(\Game_Inst.N_275_0 ),
            .ltout(\Game_Inst.N_275_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNO_0_2_LC_6_8_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNO_0_2_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNO_0_2_LC_6_8_4 .LUT_INIT=16'b0110001011101010;
    LogicCell40 \Game_Inst.r_Index_RNO_0_2_LC_6_8_4  (
            .in0(N__5958),
            .in1(N__5976),
            .in2(N__5592),
            .in3(N__5701),
            .lcout(),
            .ltout(\Game_Inst.N_268_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_2_LC_6_8_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_2_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Index_2_LC_6_8_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \Game_Inst.r_Index_2_LC_6_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5589),
            .in3(N__5584),
            .lcout(\Game_Inst.r_IndexZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8412),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_1__RNIB13I_0_LC_6_8_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_1__RNIB13I_0_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_1__RNIB13I_0_LC_6_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Game_Inst.r_Pattern_1__RNIB13I_0_LC_6_8_6  (
            .in0(N__6393),
            .in1(N__6563),
            .in2(_gnd_net_),
            .in3(N__6387),
            .lcout(),
            .ltout(\Game_Inst.r_Pattern_1__RNIB13IZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNI9R7G1_1_LC_6_8_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNI9R7G1_1_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNI9R7G1_1_LC_6_8_7 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \Game_Inst.r_Index_RNI9R7G1_1_LC_6_8_7  (
            .in0(N__6000),
            .in1(N__5957),
            .in2(N__5571),
            .in3(N__5568),
            .lcout(\Game_Inst.un1_r_Pattern_0__7_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNII65J1_1_LC_6_9_0 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNII65J1_1_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNII65J1_1_LC_6_9_0 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNII65J1_1_LC_6_9_0  (
            .in0(N__6161),
            .in1(N__5768),
            .in2(N__5898),
            .in3(N__5789),
            .lcout(\Game_Inst.SUM_i_o3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNIB3TT2_2_LC_6_9_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNIB3TT2_2_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNIB3TT2_2_LC_6_9_1 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \Game_Inst.r_Index_RNIB3TT2_2_LC_6_9_1  (
            .in0(N__5960),
            .in1(N__6519),
            .in2(N__6618),
            .in3(N__5556),
            .lcout(\Game_Inst.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNID69B_1_LC_6_9_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNID69B_1_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNID69B_1_LC_6_9_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Game_Inst.r_Index_RNID69B_1_LC_6_9_2  (
            .in0(N__6570),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6002),
            .lcout(\Game_Inst.N_276_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_5__RNIL3KJ_1_LC_6_9_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_5__RNIL3KJ_1_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_5__RNIL3KJ_1_LC_6_9_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Game_Inst.r_Pattern_5__RNIL3KJ_1_LC_6_9_3  (
            .in0(N__7212),
            .in1(N__7434),
            .in2(_gnd_net_),
            .in3(N__6569),
            .lcout(),
            .ltout(\Game_Inst.r_Pattern_5__RNIL3KJZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Index_RNIJBTT2_2_LC_6_9_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Index_RNIJBTT2_2_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Index_RNIJBTT2_2_LC_6_9_4 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \Game_Inst.r_Index_RNIJBTT2_2_LC_6_9_4  (
            .in0(N__6357),
            .in1(N__5959),
            .in2(N__5934),
            .in3(N__5931),
            .lcout(\Game_Inst.N_31 ),
            .ltout(\Game_Inst.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_ID_RNIBUVL6_0_LC_6_9_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_ID_RNIBUVL6_0_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Button_ID_RNIBUVL6_0_LC_6_9_5 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Game_Inst.r_Button_ID_RNIBUVL6_0_LC_6_9_5  (
            .in0(N__6027),
            .in1(N__6180),
            .in2(N__5925),
            .in3(N__7900),
            .lcout(\Game_Inst.un1_r_Pattern_0__1_i_0 ),
            .ltout(\Game_Inst.un1_r_Pattern_0__1_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNIVHER7_2_LC_6_9_6 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNIVHER7_2_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNIVHER7_2_LC_6_9_6 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \Game_Inst.r_SM_Main_RNIVHER7_2_LC_6_9_6  (
            .in0(N__5894),
            .in1(N__5867),
            .in2(N__5793),
            .in3(N__5790),
            .lcout(),
            .ltout(\Game_Inst.N_269_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI1KGC8_1_LC_6_9_7 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI1KGC8_1_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI1KGC8_1_LC_6_9_7 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \Game_Inst.r_SM_Main_RNI1KGC8_1_LC_6_9_7  (
            .in0(N__5769),
            .in1(_gnd_net_),
            .in2(N__5706),
            .in3(N__6162),
            .lcout(\Game_Inst.N_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_4_RNITCGR_LC_6_10_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_4_RNITCGR_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Switch_4_RNITCGR_LC_6_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Game_Inst.r_Switch_4_RNITCGR_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__7489),
            .in2(_gnd_net_),
            .in3(N__5688),
            .lcout(\Game_Inst.un1_i_Switch_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_4_LC_6_10_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_4_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Switch_4_LC_6_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Switch_4_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7490),
            .lcout(\Game_Inst.r_SwitchZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8423),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_ID_0_LC_6_10_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_ID_0_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Button_ID_0_LC_6_10_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \Game_Inst.r_Button_ID_0_LC_6_10_4  (
            .in0(N__6088),
            .in1(N__6134),
            .in2(_gnd_net_),
            .in3(N__6491),
            .lcout(\Game_Inst.r_Button_IDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8423),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main33_i_o3_LC_6_10_5 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main33_i_o3_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main33_i_o3_LC_6_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Game_Inst.r_SM_Main33_i_o3_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__7548),
            .in2(_gnd_net_),
            .in3(N__6087),
            .lcout(\Game_Inst.N_270_li ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Button_ID_1_LC_6_10_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Button_ID_1_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Button_ID_1_LC_6_10_7 .LUT_INIT=16'b1001100100001001;
    LogicCell40 \Game_Inst.r_Button_ID_1_LC_6_10_7  (
            .in0(N__6492),
            .in1(N__7358),
            .in2(N__6138),
            .in3(N__6089),
            .lcout(\Game_Inst.r_Button_IDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8423),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_1_cry_1_c_LC_6_13_0 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_1_cry_1_c_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_1_cry_1_c_LC_6_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_SW2.r_Count_1_cry_1_c_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__7695),
            .in2(N__7671),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_13_0_),
            .carryout(\Debounce_SW2.r_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_2_LC_6_13_1 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_2_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_2_LC_6_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_2_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(N__6477),
            .in2(_gnd_net_),
            .in3(N__6018),
            .lcout(\Debounce_SW2.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_1 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_2 ),
            .clk(N__8436),
            .ce(),
            .sr(N__7646));
    defparam \Debounce_SW2.r_Count_3_LC_6_13_2 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_3_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_3_LC_6_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_3_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(N__6464),
            .in2(_gnd_net_),
            .in3(N__6015),
            .lcout(\Debounce_SW2.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_2 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_3 ),
            .clk(N__8436),
            .ce(),
            .sr(N__7646));
    defparam \Debounce_SW2.r_Count_4_LC_6_13_3 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_4_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_4_LC_6_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_4_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(N__6428),
            .in2(_gnd_net_),
            .in3(N__6012),
            .lcout(\Debounce_SW2.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_3 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_4 ),
            .clk(N__8436),
            .ce(),
            .sr(N__7646));
    defparam \Debounce_SW2.r_Count_5_LC_6_13_4 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_5_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_5_LC_6_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_5_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(N__6858),
            .in2(_gnd_net_),
            .in3(N__6009),
            .lcout(\Debounce_SW2.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_4 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_5 ),
            .clk(N__8436),
            .ce(),
            .sr(N__7646));
    defparam \Debounce_SW2.r_Count_6_LC_6_13_5 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_6_LC_6_13_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_6_LC_6_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_6_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(N__6449),
            .in2(_gnd_net_),
            .in3(N__6006),
            .lcout(\Debounce_SW2.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_5 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_6 ),
            .clk(N__8436),
            .ce(),
            .sr(N__7646));
    defparam \Debounce_SW2.r_Count_7_LC_6_13_6 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_7_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_7_LC_6_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_7_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__6635),
            .in2(_gnd_net_),
            .in3(N__6207),
            .lcout(\Debounce_SW2.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_6 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_7 ),
            .clk(N__8436),
            .ce(),
            .sr(N__7646));
    defparam \Debounce_SW2.r_Count_8_LC_6_13_7 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_8_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_8_LC_6_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_8_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(N__6879),
            .in2(_gnd_net_),
            .in3(N__6204),
            .lcout(\Debounce_SW2.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_7 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_8 ),
            .clk(N__8436),
            .ce(),
            .sr(N__7646));
    defparam \Debounce_SW2.r_Count_9_LC_6_14_0 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_9_LC_6_14_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_9_LC_6_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_9_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__6828),
            .in2(_gnd_net_),
            .in3(N__6201),
            .lcout(\Debounce_SW2.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\Debounce_SW2.r_Count_1_cry_9 ),
            .clk(N__8443),
            .ce(),
            .sr(N__7645));
    defparam \Debounce_SW2.r_Count_10_LC_6_14_1 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_10_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_10_LC_6_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_10_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__6816),
            .in2(_gnd_net_),
            .in3(N__6198),
            .lcout(\Debounce_SW2.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_9 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_10 ),
            .clk(N__8443),
            .ce(),
            .sr(N__7645));
    defparam \Debounce_SW2.r_Count_11_LC_6_14_2 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_11_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_11_LC_6_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_11_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__6411),
            .in2(_gnd_net_),
            .in3(N__6195),
            .lcout(\Debounce_SW2.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_10 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_11 ),
            .clk(N__8443),
            .ce(),
            .sr(N__7645));
    defparam \Debounce_SW2.r_Count_12_LC_6_14_3 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_12_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_12_LC_6_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_12_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__7020),
            .in2(_gnd_net_),
            .in3(N__6192),
            .lcout(\Debounce_SW2.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_11 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_12 ),
            .clk(N__8443),
            .ce(),
            .sr(N__7645));
    defparam \Debounce_SW2.r_Count_13_LC_6_14_4 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_13_LC_6_14_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_13_LC_6_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_13_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__6711),
            .in2(_gnd_net_),
            .in3(N__6189),
            .lcout(\Debounce_SW2.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_12 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_13 ),
            .clk(N__8443),
            .ce(),
            .sr(N__7645));
    defparam \Debounce_SW2.r_Count_14_LC_6_14_5 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_14_LC_6_14_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_14_LC_6_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_14_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(N__6696),
            .in2(_gnd_net_),
            .in3(N__6186),
            .lcout(\Debounce_SW2.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_13 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_14 ),
            .clk(N__8443),
            .ce(),
            .sr(N__7645));
    defparam \Debounce_SW2.r_Count_15_LC_6_14_6 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_15_LC_6_14_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_15_LC_6_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_15_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(N__6726),
            .in2(_gnd_net_),
            .in3(N__6183),
            .lcout(\Debounce_SW2.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_14 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_15 ),
            .clk(N__8443),
            .ce(),
            .sr(N__7645));
    defparam \Debounce_SW2.r_Count_16_LC_6_14_7 .C_ON=1'b1;
    defparam \Debounce_SW2.r_Count_16_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_16_LC_6_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW2.r_Count_16_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(N__6671),
            .in2(_gnd_net_),
            .in3(N__6276),
            .lcout(\Debounce_SW2.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_SW2.r_Count_1_cry_15 ),
            .carryout(\Debounce_SW2.r_Count_1_cry_16 ),
            .clk(N__8443),
            .ce(),
            .sr(N__7645));
    defparam \Debounce_SW2.r_Count_17_LC_6_15_0 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_17_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_17_LC_6_15_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_SW2.r_Count_17_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(N__6654),
            .in2(_gnd_net_),
            .in3(N__6273),
            .lcout(\Debounce_SW2.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8446),
            .ce(),
            .sr(N__7644));
    defparam \Debounce_SW4.r_State_RNI9SDT2_LC_7_4_4 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_RNI9SDT2_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_State_RNI9SDT2_LC_7_4_4 .LUT_INIT=16'b1010010111101101;
    LogicCell40 \Debounce_SW4.r_State_RNI9SDT2_LC_7_4_4  (
            .in0(N__7476),
            .in1(N__6333),
            .in2(N__6257),
            .in3(N__6213),
            .lcout(\Debounce_SW4.r_Count12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_State_RNO_1_LC_7_5_0 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_RNO_1_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_State_RNO_1_LC_7_5_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Debounce_SW4.r_State_RNO_1_LC_7_5_0  (
            .in0(N__6996),
            .in1(N__7142),
            .in2(N__6324),
            .in3(N__7164),
            .lcout(\Debounce_SW4.r_Count13_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_State_RNO_0_LC_7_5_2 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_RNO_0_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_State_RNO_0_LC_7_5_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Debounce_SW4.r_State_RNO_0_LC_7_5_2  (
            .in0(N__7181),
            .in1(N__6225),
            .in2(N__6900),
            .in3(N__6315),
            .lcout(),
            .ltout(\Debounce_SW4.r_Count13_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_State_LC_7_5_3 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_State_LC_7_5_3 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Debounce_SW4.r_State_LC_7_5_3  (
            .in0(N__6261),
            .in1(N__6234),
            .in2(N__6228),
            .in3(N__7477),
            .lcout(w_Switch_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8431),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNID2KD_4_LC_7_5_4 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNID2KD_4_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNID2KD_4_LC_7_5_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Debounce_SW4.r_Count_RNID2KD_4_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__6914),
            .in2(_gnd_net_),
            .in3(N__6929),
            .lcout(\Debounce_SW4.r_Count13_1 ),
            .ltout(\Debounce_SW4.r_Count13_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNIC1GM1_6_LC_7_5_5 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNIC1GM1_6_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNIC1GM1_6_LC_7_5_5 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \Debounce_SW4.r_Count_RNIC1GM1_6_LC_7_5_5  (
            .in0(N__7201),
            .in1(N__6895),
            .in2(N__6219),
            .in3(N__6995),
            .lcout(),
            .ltout(\Debounce_SW4.un1_r_Count_8lt11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNIJ6T62_12_LC_7_5_6 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNIJ6T62_12_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNIJ6T62_12_LC_7_5_6 .LUT_INIT=16'b0001001100010001;
    LogicCell40 \Debounce_SW4.r_Count_RNIJ6T62_12_LC_7_5_6  (
            .in0(N__7099),
            .in1(N__7079),
            .in2(N__6216),
            .in3(N__6339),
            .lcout(\Debounce_SW4.un1_r_Count_8lt17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNISL0F_10_LC_7_5_7 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNISL0F_10_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNISL0F_10_LC_7_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Debounce_SW4.r_Count_RNISL0F_10_LC_7_5_7  (
            .in0(N__7141),
            .in1(N__7162),
            .in2(N__7125),
            .in3(N__7180),
            .lcout(\Debounce_SW4.un1_r_Count_8lto11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_RNI2BP2_17_LC_7_6_0 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNI2BP2_17_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNI2BP2_17_LC_7_6_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW4.r_Count_RNI2BP2_17_LC_7_6_0  (
            .in0(N__7309),
            .in1(N__7033),
            .in2(N__7289),
            .in3(N__7051),
            .lcout(\Debounce_SW4.un1_r_Count_8lto17_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_State_RNO_3_LC_7_6_5 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_RNO_3_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_State_RNO_3_LC_7_6_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Debounce_SW4.r_State_RNO_3_LC_7_6_5  (
            .in0(N__7100),
            .in1(N__7123),
            .in2(N__7080),
            .in3(N__7202),
            .lcout(\Debounce_SW4.r_Count13_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_State_RNO_2_LC_7_6_6 .C_ON=1'b0;
    defparam \Debounce_SW4.r_State_RNO_2_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_State_RNO_2_LC_7_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW4.r_State_RNO_2_LC_7_6_6  (
            .in0(N__7310),
            .in1(N__7034),
            .in2(N__7290),
            .in3(N__7052),
            .lcout(\Debounce_SW4.r_Count13_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_1__RNID33I_1_LC_7_7_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_1__RNID33I_1_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_1__RNID33I_1_LC_7_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Game_Inst.r_Pattern_1__RNID33I_1_LC_7_7_1  (
            .in0(N__6294),
            .in1(N__6564),
            .in2(_gnd_net_),
            .in3(N__6399),
            .lcout(\Game_Inst.r_Pattern_1__RNID33IZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_2__RNIHJRI_1_LC_7_7_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_2__RNIHJRI_1_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_2__RNIHJRI_1_LC_7_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Game_Inst.r_Pattern_2__RNIHJRI_1_LC_7_7_2  (
            .in0(N__6565),
            .in1(N__6288),
            .in2(_gnd_net_),
            .in3(N__6282),
            .lcout(\Game_Inst.r_Pattern_2__RNIHJRIZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_0__1_LC_7_7_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_0__1_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_0__1_LC_7_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_0__1_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6609),
            .lcout(\Game_Inst.r_Pattern_0_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8424),
            .ce(N__7401),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_2__1_LC_7_7_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_2__1_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_2__1_LC_7_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_2__1_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7257),
            .lcout(\Game_Inst.r_Pattern_2_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8424),
            .ce(N__7401),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_3__1_LC_7_8_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_3__1_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_3__1_LC_7_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_3__1_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7269),
            .lcout(\Game_Inst.r_Pattern_3_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8417),
            .ce(N__7400),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_1__1_LC_7_8_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_1__1_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_1__1_LC_7_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_1__1_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6369),
            .lcout(\Game_Inst.r_Pattern_1_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8417),
            .ce(N__7400),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_0__0_LC_7_8_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_0__0_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_0__0_LC_7_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_0__0_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7716),
            .lcout(\Game_Inst.r_Pattern_0_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8417),
            .ce(N__7400),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_1__0_LC_7_8_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_1__0_LC_7_8_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_1__0_LC_7_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_1__0_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6594),
            .lcout(\Game_Inst.r_Pattern_1_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8417),
            .ce(N__7400),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_2__0_LC_7_8_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_2__0_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_2__0_LC_7_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_2__0_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6351),
            .lcout(\Game_Inst.r_Pattern_2_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8417),
            .ce(N__7400),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_3__0_LC_7_8_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_3__0_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_3__0_LC_7_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_3__0_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7242),
            .lcout(\Game_Inst.r_Pattern_3_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8417),
            .ce(N__7400),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_4_LC_7_9_0 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_4_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_4_LC_7_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_4_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6368),
            .lcout(\Game_Inst.w_LFSR_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8425),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_3_LC_7_9_1 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_3_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_3_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_3_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6593),
            .lcout(\Game_Inst.w_LFSR_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8425),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_6__RNIPJCK_1_LC_7_9_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_6__RNIPJCK_1_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_6__RNIPJCK_1_LC_7_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Game_Inst.r_Pattern_6__RNIPJCK_1_LC_7_9_2  (
            .in0(N__6568),
            .in1(N__7407),
            .in2(_gnd_net_),
            .in3(N__7419),
            .lcout(\Game_Inst.r_Pattern_6__RNIPJCKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_1_LC_7_9_3 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_1_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_1_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_1_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7715),
            .lcout(\Game_Inst.w_LFSR_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8425),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_5_LC_7_9_4 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_5_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_5_LC_7_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_5_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6350),
            .lcout(\Game_Inst.w_LFSR_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8425),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_6__RNINHCK_0_LC_7_9_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_6__RNINHCK_0_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_6__RNINHCK_0_LC_7_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Game_Inst.r_Pattern_6__RNINHCK_0_LC_7_9_5  (
            .in0(N__7413),
            .in1(N__7425),
            .in2(_gnd_net_),
            .in3(N__6567),
            .lcout(\Game_Inst.r_Pattern_6__RNINHCKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_2_LC_7_9_6 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_2_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_2_LC_7_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_2_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6605),
            .lcout(\Game_Inst.w_LFSR_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8425),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_5__RNIJ1KJ_0_LC_7_9_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_5__RNIJ1KJ_0_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Pattern_5__RNIJ1KJ_0_LC_7_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Game_Inst.r_Pattern_5__RNIJ1KJ_0_LC_7_9_7  (
            .in0(N__7440),
            .in1(N__7218),
            .in2(_gnd_net_),
            .in3(N__6566),
            .lcout(\Game_Inst.r_Pattern_5__RNIJ1KJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_2_RNIABK13_LC_7_10_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_2_RNIABK13_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Switch_2_RNIABK13_LC_7_10_4 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \Game_Inst.r_Switch_2_RNIABK13_LC_7_10_4  (
            .in0(N__7348),
            .in1(N__7332),
            .in2(N__6509),
            .in3(N__7566),
            .lcout(\Game_Inst.r_Button_ID_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_LC_7_11_3 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_State_LC_7_11_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \Debounce_SW2.r_State_LC_7_11_3  (
            .in0(N__6483),
            .in1(N__6843),
            .in2(N__6770),
            .in3(N__7567),
            .lcout(w_Switch_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8430),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_RNO_0_LC_7_12_2 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_RNO_0_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_State_RNO_0_LC_7_12_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Debounce_SW2.r_State_RNO_0_LC_7_12_2  (
            .in0(N__6450),
            .in1(N__6429),
            .in2(N__6804),
            .in3(N__6792),
            .lcout(\Debounce_SW2.r_Count13_0_a7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNI60D51_1_LC_7_13_1 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNI60D51_1_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNI60D51_1_LC_7_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW2.r_Count_RNI60D51_1_LC_7_13_1  (
            .in0(N__6476),
            .in1(N__7663),
            .in2(N__6465),
            .in3(N__7689),
            .lcout(\Debounce_SW2.r_Count13_10 ),
            .ltout(\Debounce_SW2.r_Count13_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNI53F12_4_LC_7_13_2 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNI53F12_4_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNI53F12_4_LC_7_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Debounce_SW2.r_Count_RNI53F12_4_LC_7_13_2  (
            .in0(N__6448),
            .in1(N__6856),
            .in2(N__6432),
            .in3(N__6427),
            .lcout(\Debounce_SW2.N_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNIQSSD_11_LC_7_13_3 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNIQSSD_11_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNIQSSD_11_LC_7_13_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Debounce_SW2.r_Count_RNIQSSD_11_LC_7_13_3  (
            .in0(N__6410),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6878),
            .lcout(\Debounce_SW2.N_23_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_RNO_1_LC_7_13_6 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_RNO_1_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_State_RNO_1_LC_7_13_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Debounce_SW2.r_State_RNO_1_LC_7_13_6  (
            .in0(N__7002),
            .in1(N__6834),
            .in2(N__6867),
            .in3(N__6857),
            .lcout(\Debounce_SW2.r_Count13_0_a7_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_RNO_2_LC_7_14_0 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_RNO_2_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_State_RNO_2_LC_7_14_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Debounce_SW2.r_State_RNO_2_LC_7_14_0  (
            .in0(N__6725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6695),
            .lcout(\Debounce_SW2.r_Count13_0_a7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNIUCEI_10_LC_7_14_1 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNIUCEI_10_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNIUCEI_10_LC_7_14_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Debounce_SW2.r_Count_RNIUCEI_10_LC_7_14_1  (
            .in0(N__6710),
            .in1(N__6827),
            .in2(_gnd_net_),
            .in3(N__6815),
            .lcout(\Debounce_SW2.N_23_2 ),
            .ltout(\Debounce_SW2.N_23_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNIKQ5B3_7_LC_7_14_2 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNIKQ5B3_7_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNIKQ5B3_7_LC_7_14_2 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \Debounce_SW2.r_Count_RNIKQ5B3_7_LC_7_14_2  (
            .in0(N__6631),
            .in1(N__6791),
            .in2(N__6780),
            .in3(N__6777),
            .lcout(),
            .ltout(\Debounce_SW2.N_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_RNI5LPJ4_LC_7_14_3 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_RNI5LPJ4_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_State_RNI5LPJ4_LC_7_14_3 .LUT_INIT=16'b1010101101010111;
    LogicCell40 \Debounce_SW2.r_State_RNI5LPJ4_LC_7_14_3  (
            .in0(N__6771),
            .in1(N__6678),
            .in2(N__6741),
            .in3(N__7577),
            .lcout(\Debounce_SW2.r_Count12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNIK46I_12_LC_7_14_4 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNIK46I_12_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNIK46I_12_LC_7_14_4 .LUT_INIT=16'b0101111101111111;
    LogicCell40 \Debounce_SW2.r_Count_RNIK46I_12_LC_7_14_4  (
            .in0(N__6724),
            .in1(N__6709),
            .in2(N__6672),
            .in3(N__7018),
            .lcout(),
            .ltout(\Debounce_SW2.un1_r_Count_8lto17_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_RNI1A9R_17_LC_7_14_5 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_RNI1A9R_17_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_Count_RNI1A9R_17_LC_7_14_5 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \Debounce_SW2.r_Count_RNI1A9R_17_LC_7_14_5  (
            .in0(N__6694),
            .in1(_gnd_net_),
            .in2(N__6681),
            .in3(N__6652),
            .lcout(\Debounce_SW2.un1_r_Count_8lto17_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_State_RNO_3_LC_7_14_6 .C_ON=1'b0;
    defparam \Debounce_SW2.r_State_RNO_3_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW2.r_State_RNO_3_LC_7_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW2.r_State_RNO_3_LC_7_14_6  (
            .in0(N__6670),
            .in1(N__6653),
            .in2(N__6636),
            .in3(N__7019),
            .lcout(\Debounce_SW2.r_Count13_0_a7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_1_LC_8_3_6 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_1_LC_8_3_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_1_LC_8_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \Debounce_SW4.r_Count_1_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(N__6983),
            .in2(_gnd_net_),
            .in3(N__7629),
            .lcout(\Debounce_SW4.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8448),
            .ce(),
            .sr(N__7601));
    defparam \Debounce_SW4.r_Count_RNIEO7R_1_LC_8_4_6 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_RNIEO7R_1_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_RNIEO7R_1_LC_8_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW4.r_Count_RNIEO7R_1_LC_8_4_6  (
            .in0(N__6962),
            .in1(N__6979),
            .in2(N__6948),
            .in3(N__7626),
            .lcout(\Debounce_SW4.r_Count13_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_1_cry_1_c_LC_8_5_0 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_1_cry_1_c_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW4.r_Count_1_cry_1_c_LC_8_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_SW4.r_Count_1_cry_1_c_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__7627),
            .in2(N__6987),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\Debounce_SW4.r_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW4.r_Count_2_LC_8_5_1 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_2_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_2_LC_8_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_2_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(N__6963),
            .in2(_gnd_net_),
            .in3(N__6951),
            .lcout(\Debounce_SW4.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_1 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_2 ),
            .clk(N__8438),
            .ce(),
            .sr(N__7602));
    defparam \Debounce_SW4.r_Count_3_LC_8_5_2 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_3_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_3_LC_8_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_3_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__6947),
            .in2(_gnd_net_),
            .in3(N__6933),
            .lcout(\Debounce_SW4.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_2 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_3 ),
            .clk(N__8438),
            .ce(),
            .sr(N__7602));
    defparam \Debounce_SW4.r_Count_4_LC_8_5_3 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_4_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_4_LC_8_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_4_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__6930),
            .in2(_gnd_net_),
            .in3(N__6918),
            .lcout(\Debounce_SW4.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_3 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_4 ),
            .clk(N__8438),
            .ce(),
            .sr(N__7602));
    defparam \Debounce_SW4.r_Count_5_LC_8_5_4 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_5_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_5_LC_8_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_5_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(N__6915),
            .in2(_gnd_net_),
            .in3(N__6903),
            .lcout(\Debounce_SW4.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_4 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_5 ),
            .clk(N__8438),
            .ce(),
            .sr(N__7602));
    defparam \Debounce_SW4.r_Count_6_LC_8_5_5 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_6_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_6_LC_8_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_6_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(N__6899),
            .in2(_gnd_net_),
            .in3(N__6882),
            .lcout(\Debounce_SW4.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_5 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_6 ),
            .clk(N__8438),
            .ce(),
            .sr(N__7602));
    defparam \Debounce_SW4.r_Count_7_LC_8_5_6 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_7_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_7_LC_8_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_7_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(N__7203),
            .in2(_gnd_net_),
            .in3(N__7185),
            .lcout(\Debounce_SW4.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_6 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_7 ),
            .clk(N__8438),
            .ce(),
            .sr(N__7602));
    defparam \Debounce_SW4.r_Count_8_LC_8_5_7 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_8_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_8_LC_8_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_8_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(N__7182),
            .in2(_gnd_net_),
            .in3(N__7167),
            .lcout(\Debounce_SW4.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_7 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_8 ),
            .clk(N__8438),
            .ce(),
            .sr(N__7602));
    defparam \Debounce_SW4.r_Count_9_LC_8_6_0 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_9_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_9_LC_8_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_9_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__7163),
            .in2(_gnd_net_),
            .in3(N__7146),
            .lcout(\Debounce_SW4.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\Debounce_SW4.r_Count_1_cry_9 ),
            .clk(N__8433),
            .ce(),
            .sr(N__7604));
    defparam \Debounce_SW4.r_Count_10_LC_8_6_1 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_10_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_10_LC_8_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_10_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__7143),
            .in2(_gnd_net_),
            .in3(N__7128),
            .lcout(\Debounce_SW4.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_9 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_10 ),
            .clk(N__8433),
            .ce(),
            .sr(N__7604));
    defparam \Debounce_SW4.r_Count_11_LC_8_6_2 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_11_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_11_LC_8_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_11_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__7124),
            .in2(_gnd_net_),
            .in3(N__7104),
            .lcout(\Debounce_SW4.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_10 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_11 ),
            .clk(N__8433),
            .ce(),
            .sr(N__7604));
    defparam \Debounce_SW4.r_Count_12_LC_8_6_3 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_12_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_12_LC_8_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_12_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__7101),
            .in2(_gnd_net_),
            .in3(N__7083),
            .lcout(\Debounce_SW4.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_11 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_12 ),
            .clk(N__8433),
            .ce(),
            .sr(N__7604));
    defparam \Debounce_SW4.r_Count_13_LC_8_6_4 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_13_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_13_LC_8_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_13_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__7078),
            .in2(_gnd_net_),
            .in3(N__7056),
            .lcout(\Debounce_SW4.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_12 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_13 ),
            .clk(N__8433),
            .ce(),
            .sr(N__7604));
    defparam \Debounce_SW4.r_Count_14_LC_8_6_5 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_14_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_14_LC_8_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_14_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__7053),
            .in2(_gnd_net_),
            .in3(N__7038),
            .lcout(\Debounce_SW4.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_13 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_14 ),
            .clk(N__8433),
            .ce(),
            .sr(N__7604));
    defparam \Debounce_SW4.r_Count_15_LC_8_6_6 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_15_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_15_LC_8_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_15_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__7035),
            .in2(_gnd_net_),
            .in3(N__7314),
            .lcout(\Debounce_SW4.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_14 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_15 ),
            .clk(N__8433),
            .ce(),
            .sr(N__7604));
    defparam \Debounce_SW4.r_Count_16_LC_8_6_7 .C_ON=1'b1;
    defparam \Debounce_SW4.r_Count_16_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_16_LC_8_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW4.r_Count_16_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__7311),
            .in2(_gnd_net_),
            .in3(N__7296),
            .lcout(\Debounce_SW4.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_SW4.r_Count_1_cry_15 ),
            .carryout(\Debounce_SW4.r_Count_1_cry_16 ),
            .clk(N__8433),
            .ce(),
            .sr(N__7604));
    defparam \Debounce_SW4.r_Count_17_LC_8_7_0 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_17_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_17_LC_8_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_SW4.r_Count_17_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__7288),
            .in2(_gnd_net_),
            .in3(N__7293),
            .lcout(\Debounce_SW4.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8427),
            .ce(),
            .sr(N__7605));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_8_LC_8_8_0 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_8_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_8_LC_8_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_8_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7268),
            .lcout(\Game_Inst.w_LFSR_Data_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8420),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_7_LC_8_8_2 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_7_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_7_LC_8_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_7_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7241),
            .lcout(\Game_Inst.w_LFSR_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8420),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_6_LC_8_8_6 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_6_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_6_LC_8_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_6_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7256),
            .lcout(\Game_Inst.w_LFSR_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8420),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_9_LC_8_8_7 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_9_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_9_LC_8_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_9_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7229),
            .lcout(\Game_Inst.w_LFSR_Data_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8420),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_4__0_LC_8_9_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_4__0_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_4__0_LC_8_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_4__0_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7230),
            .lcout(\Game_Inst.r_Pattern_4_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8428),
            .ce(N__7393),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_4__1_LC_8_9_1 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_4__1_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_4__1_LC_8_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_4__1_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7826),
            .lcout(\Game_Inst.r_Pattern_4_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8428),
            .ce(N__7393),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_5__0_LC_8_9_2 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_5__0_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_5__0_LC_8_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_5__0_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7815),
            .lcout(\Game_Inst.r_Pattern_5_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8428),
            .ce(N__7393),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_5__1_LC_8_9_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_5__1_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_5__1_LC_8_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_5__1_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7779),
            .lcout(\Game_Inst.r_Pattern_5_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8428),
            .ce(N__7393),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_6__0_LC_8_9_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_6__0_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_6__0_LC_8_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_6__0_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7767),
            .lcout(\Game_Inst.r_Pattern_6_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8428),
            .ce(N__7393),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_6__1_LC_8_9_5 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_6__1_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_6__1_LC_8_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_6__1_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7803),
            .lcout(\Game_Inst.r_Pattern_6_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8428),
            .ce(N__7393),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_7__0_LC_8_9_6 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_7__0_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_7__0_LC_8_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.r_Pattern_7__0_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7791),
            .lcout(\Game_Inst.r_Pattern_7_Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8428),
            .ce(N__7393),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Pattern_7__1_LC_8_9_7 .C_ON=1'b0;
    defparam \Game_Inst.r_Pattern_7__1_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Pattern_7__1_LC_8_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Game_Inst.r_Pattern_7__1_LC_8_9_7  (
            .in0(N__7755),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.r_Pattern_7_Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8428),
            .ce(N__7393),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_3_RNIK1CC1_LC_8_10_0 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_3_RNIK1CC1_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_Switch_3_RNIK1CC1_LC_8_10_0 .LUT_INIT=16'b1111010100110001;
    LogicCell40 \Game_Inst.r_Switch_3_RNIK1CC1_LC_8_10_0  (
            .in0(N__7320),
            .in1(N__7331),
            .in2(N__8489),
            .in3(N__7555),
            .lcout(\Game_Inst.r_Button_ID_2_sm0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_2_LC_8_10_3 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_2_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Switch_2_LC_8_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Game_Inst.r_Switch_2_LC_8_10_3  (
            .in0(N__7556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.r_SwitchZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8432),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_Switch_3_LC_8_10_4 .C_ON=1'b0;
    defparam \Game_Inst.r_Switch_3_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.r_Switch_3_LC_8_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Game_Inst.r_Switch_3_LC_8_10_4  (
            .in0(N__8485),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Game_Inst.r_SwitchZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8432),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_19_LC_8_11_0 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_19_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_19_LC_8_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_19_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7968),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8437),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_21_LC_8_11_2 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_21_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_21_LC_8_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_21_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7725),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8437),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_20_LC_8_11_4 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_20_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_20_LC_8_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_20_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7737),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8437),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_0_LC_8_11_6 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_0_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_0_LC_8_11_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_0_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__7731),
            .in2(_gnd_net_),
            .in3(N__7724),
            .lcout(\Game_Inst.w_LFSR_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8437),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW2.r_Count_0_LC_8_13_2 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_0_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_0_LC_8_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_SW2.r_Count_0_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7693),
            .lcout(\Debounce_SW2.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8447),
            .ce(),
            .sr(N__7647));
    defparam \Debounce_SW2.r_Count_1_LC_8_13_5 .C_ON=1'b0;
    defparam \Debounce_SW2.r_Count_1_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW2.r_Count_1_LC_8_13_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Debounce_SW2.r_Count_1_LC_8_13_5  (
            .in0(N__7694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7667),
            .lcout(\Debounce_SW2.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8447),
            .ce(),
            .sr(N__7647));
    defparam \Debounce_SW4.r_Count_0_LC_9_4_6 .C_ON=1'b0;
    defparam \Debounce_SW4.r_Count_0_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW4.r_Count_0_LC_9_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_SW4.r_Count_0_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7628),
            .lcout(\Debounce_SW4.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8449),
            .ce(),
            .sr(N__7603));
    defparam \Game_Inst.r_SM_Main_RNI776H6_1_LC_9_7_1 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI776H6_1_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI776H6_1_LC_9_7_1 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \Game_Inst.r_SM_Main_RNI776H6_1_LC_9_7_1  (
            .in0(N__7915),
            .in1(N__7882),
            .in2(N__7856),
            .in3(N__7582),
            .lcout(Game_Inst_o_LED_2_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI9NUI6_1_LC_9_7_2 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI9NUI6_1_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI9NUI6_1_LC_9_7_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Game_Inst.r_SM_Main_RNI9NUI6_1_LC_9_7_2  (
            .in0(N__7884),
            .in1(N__7855),
            .in2(N__7494),
            .in3(N__7917),
            .lcout(Game_Inst_o_LED_4_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.r_SM_Main_RNI8F2A6_1_LC_9_7_3 .C_ON=1'b0;
    defparam \Game_Inst.r_SM_Main_RNI8F2A6_1_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \Game_Inst.r_SM_Main_RNI8F2A6_1_LC_9_7_3 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \Game_Inst.r_SM_Main_RNI8F2A6_1_LC_9_7_3  (
            .in0(N__7916),
            .in1(N__7883),
            .in2(N__7857),
            .in3(N__8490),
            .lcout(Game_Inst_o_LED_3_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_10_LC_9_9_1 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_10_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_10_LC_9_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_10_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7827),
            .lcout(\Game_Inst.w_LFSR_Data_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8434),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_11_LC_9_9_2 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_11_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_11_LC_9_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_11_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7814),
            .lcout(\Game_Inst.w_LFSR_Data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8434),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_15_LC_9_9_3 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_15_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_15_LC_9_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_15_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7790),
            .lcout(\Game_Inst.w_LFSR_Data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8434),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_13_LC_9_9_4 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_13_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_13_LC_9_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_13_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7766),
            .lcout(\Game_Inst.w_LFSR_Data_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8434),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_14_LC_9_9_5 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_14_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_14_LC_9_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_14_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7802),
            .lcout(\Game_Inst.w_LFSR_Data_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8434),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_12_LC_9_9_7 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_12_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_12_LC_9_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_12_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7778),
            .lcout(\Game_Inst.w_LFSR_Data_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8434),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_17_LC_9_10_1 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_17_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_17_LC_9_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_17_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7743),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8439),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_16_LC_9_10_4 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_16_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_16_LC_9_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_16_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7754),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8439),
            .ce(),
            .sr(_gnd_net_));
    defparam \Game_Inst.LFSR_Inst.r_LFSR_18_LC_9_10_7 .C_ON=1'b0;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_18_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \Game_Inst.LFSR_Inst.r_LFSR_18_LC_9_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Game_Inst.LFSR_Inst.r_LFSR_18_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7974),
            .lcout(\Game_Inst.LFSR_Inst.r_LFSRZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8439),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_RNO_0_LC_11_8_0 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_RNO_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_State_RNO_0_LC_11_8_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Debounce_SW3.r_State_RNO_0_LC_11_8_0  (
            .in0(N__8084),
            .in1(N__8063),
            .in2(N__7959),
            .in3(N__7950),
            .lcout(\Debounce_SW3.r_Count13_0_a7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNIACA_1_LC_11_8_2 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNIACA_1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNIACA_1_LC_11_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW3.r_Count_RNIACA_1_LC_11_8_2  (
            .in0(N__7931),
            .in1(N__8170),
            .in2(N__8103),
            .in3(N__8151),
            .lcout(\Debounce_SW3.r_Count13_10 ),
            .ltout(\Debounce_SW3.r_Count13_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNICGI_4_LC_11_8_3 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNICGI_4_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNICGI_4_LC_11_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Debounce_SW3.r_Count_RNICGI_4_LC_11_8_3  (
            .in0(N__8062),
            .in1(N__8539),
            .in2(N__7962),
            .in3(N__8083),
            .lcout(\Debounce_SW3.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNISJM2_8_LC_11_8_4 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNISJM2_8_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNISJM2_8_LC_11_8_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Debounce_SW3.r_Count_RNISJM2_8_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__7992),
            .in2(_gnd_net_),
            .in3(N__8042),
            .lcout(\Debounce_SW3.N_18_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNI1GA5_9_LC_11_8_5 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNI1GA5_9_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNI1GA5_9_LC_11_8_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Debounce_SW3.r_Count_RNI1GA5_9_LC_11_8_5  (
            .in0(N__8010),
            .in1(N__8028),
            .in2(_gnd_net_),
            .in3(N__8286),
            .lcout(\Debounce_SW3.N_18_2 ),
            .ltout(\Debounce_SW3.N_18_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNI1DM8_7_LC_11_8_6 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNI1DM8_7_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNI1DM8_7_LC_11_8_6 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \Debounce_SW3.r_Count_RNI1DM8_7_LC_11_8_6  (
            .in0(N__8578),
            .in1(N__7949),
            .in2(N__7941),
            .in3(N__7938),
            .lcout(\Debounce_SW3.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_1_cry_1_c_LC_11_9_0 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_1_cry_1_c_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_1_cry_1_c_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Debounce_SW3.r_Count_1_cry_1_c_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__8152),
            .in2(N__8175),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\Debounce_SW3.r_Count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_2_LC_11_9_1 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_2_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_2_LC_11_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_2_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__7932),
            .in2(_gnd_net_),
            .in3(N__7920),
            .lcout(\Debounce_SW3.r_CountZ0Z_2 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_1 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_2 ),
            .clk(N__8441),
            .ce(),
            .sr(N__8130));
    defparam \Debounce_SW3.r_Count_3_LC_11_9_2 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_3_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_3_LC_11_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_3_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__8102),
            .in2(_gnd_net_),
            .in3(N__8088),
            .lcout(\Debounce_SW3.r_CountZ0Z_3 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_2 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_3 ),
            .clk(N__8441),
            .ce(),
            .sr(N__8130));
    defparam \Debounce_SW3.r_Count_4_LC_11_9_3 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_4_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_4_LC_11_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_4_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__8085),
            .in2(_gnd_net_),
            .in3(N__8070),
            .lcout(\Debounce_SW3.r_CountZ0Z_4 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_3 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_4 ),
            .clk(N__8441),
            .ce(),
            .sr(N__8130));
    defparam \Debounce_SW3.r_Count_5_LC_11_9_4 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_5_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_5_LC_11_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_5_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__8540),
            .in2(_gnd_net_),
            .in3(N__8067),
            .lcout(\Debounce_SW3.r_CountZ0Z_5 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_4 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_5 ),
            .clk(N__8441),
            .ce(),
            .sr(N__8130));
    defparam \Debounce_SW3.r_Count_6_LC_11_9_5 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_6_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_6_LC_11_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_6_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__8064),
            .in2(_gnd_net_),
            .in3(N__8049),
            .lcout(\Debounce_SW3.r_CountZ0Z_6 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_5 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_6 ),
            .clk(N__8441),
            .ce(),
            .sr(N__8130));
    defparam \Debounce_SW3.r_Count_7_LC_11_9_6 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_7_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_7_LC_11_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_7_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__8582),
            .in2(_gnd_net_),
            .in3(N__8046),
            .lcout(\Debounce_SW3.r_CountZ0Z_7 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_6 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_7 ),
            .clk(N__8441),
            .ce(),
            .sr(N__8130));
    defparam \Debounce_SW3.r_Count_8_LC_11_9_7 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_8_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_8_LC_11_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_8_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__8043),
            .in2(_gnd_net_),
            .in3(N__8031),
            .lcout(\Debounce_SW3.r_CountZ0Z_8 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_7 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_8 ),
            .clk(N__8441),
            .ce(),
            .sr(N__8130));
    defparam \Debounce_SW3.r_Count_9_LC_11_10_0 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_9_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_9_LC_11_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_9_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__8027),
            .in2(_gnd_net_),
            .in3(N__8013),
            .lcout(\Debounce_SW3.r_CountZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\Debounce_SW3.r_Count_1_cry_9 ),
            .clk(N__8444),
            .ce(),
            .sr(N__8132));
    defparam \Debounce_SW3.r_Count_10_LC_11_10_1 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_10_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_10_LC_11_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_10_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__8009),
            .in2(_gnd_net_),
            .in3(N__7995),
            .lcout(\Debounce_SW3.r_CountZ0Z_10 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_9 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_10 ),
            .clk(N__8444),
            .ce(),
            .sr(N__8132));
    defparam \Debounce_SW3.r_Count_11_LC_11_10_2 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_11_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_11_LC_11_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_11_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__7991),
            .in2(_gnd_net_),
            .in3(N__7977),
            .lcout(\Debounce_SW3.r_CountZ0Z_11 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_10 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_11 ),
            .clk(N__8444),
            .ce(),
            .sr(N__8132));
    defparam \Debounce_SW3.r_Count_12_LC_11_10_3 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_12_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_12_LC_11_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_12_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__8247),
            .in2(_gnd_net_),
            .in3(N__8193),
            .lcout(\Debounce_SW3.r_CountZ0Z_12 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_11 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_12 ),
            .clk(N__8444),
            .ce(),
            .sr(N__8132));
    defparam \Debounce_SW3.r_Count_13_LC_11_10_4 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_13_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_13_LC_11_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_13_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__8285),
            .in2(_gnd_net_),
            .in3(N__8190),
            .lcout(\Debounce_SW3.r_CountZ0Z_13 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_12 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_13 ),
            .clk(N__8444),
            .ce(),
            .sr(N__8132));
    defparam \Debounce_SW3.r_Count_14_LC_11_10_5 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_14_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_14_LC_11_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_14_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__8214),
            .in2(_gnd_net_),
            .in3(N__8187),
            .lcout(\Debounce_SW3.r_CountZ0Z_14 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_13 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_14 ),
            .clk(N__8444),
            .ce(),
            .sr(N__8132));
    defparam \Debounce_SW3.r_Count_15_LC_11_10_6 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_15_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_15_LC_11_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_15_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__8301),
            .in2(_gnd_net_),
            .in3(N__8184),
            .lcout(\Debounce_SW3.r_CountZ0Z_15 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_14 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_15 ),
            .clk(N__8444),
            .ce(),
            .sr(N__8132));
    defparam \Debounce_SW3.r_Count_16_LC_11_10_7 .C_ON=1'b1;
    defparam \Debounce_SW3.r_Count_16_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_16_LC_11_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Debounce_SW3.r_Count_16_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__8264),
            .in2(_gnd_net_),
            .in3(N__8181),
            .lcout(\Debounce_SW3.r_CountZ0Z_16 ),
            .ltout(),
            .carryin(\Debounce_SW3.r_Count_1_cry_15 ),
            .carryout(\Debounce_SW3.r_Count_1_cry_16 ),
            .clk(N__8444),
            .ce(),
            .sr(N__8132));
    defparam \Debounce_SW3.r_Count_17_LC_11_11_0 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_17_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_17_LC_11_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Debounce_SW3.r_Count_17_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__8232),
            .in2(_gnd_net_),
            .in3(N__8178),
            .lcout(\Debounce_SW3.r_CountZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8450),
            .ce(),
            .sr(N__8133));
    defparam \Debounce_SW3.r_Count_1_LC_12_8_0 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_1_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_1_LC_12_8_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \Debounce_SW3.r_Count_1_LC_12_8_0  (
            .in0(N__8154),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8174),
            .lcout(\Debounce_SW3.r_CountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8440),
            .ce(),
            .sr(N__8131));
    defparam \Debounce_SW3.r_Count_0_LC_12_8_5 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_0_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_Count_0_LC_12_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Debounce_SW3.r_Count_0_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8153),
            .lcout(\Debounce_SW3.r_CountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8440),
            .ce(),
            .sr(N__8131));
    defparam \Debounce_SW3.r_State_RNIQSU81_LC_12_9_3 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_RNIQSU81_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_State_RNIQSU81_LC_12_9_3 .LUT_INIT=16'b1010010110110111;
    LogicCell40 \Debounce_SW3.r_State_RNIQSU81_LC_12_9_3  (
            .in0(N__8477),
            .in1(N__8199),
            .in2(N__8523),
            .in3(N__8115),
            .lcout(\Debounce_SW3.r_Count12_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_RNO_2_LC_12_10_1 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_RNO_2_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_State_RNO_2_LC_12_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Debounce_SW3.r_State_RNO_2_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__8213),
            .in2(_gnd_net_),
            .in3(N__8300),
            .lcout(\Debounce_SW3.r_Count13_0_a7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_RNO_3_LC_12_10_3 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_RNO_3_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_State_RNO_3_LC_12_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Debounce_SW3.r_State_RNO_3_LC_12_10_3  (
            .in0(N__8246),
            .in1(N__8231),
            .in2(N__8583),
            .in3(N__8263),
            .lcout(),
            .ltout(\Debounce_SW3.r_Count13_0_a7_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_RNO_1_LC_12_10_4 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_RNO_1_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_State_RNO_1_LC_12_10_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Debounce_SW3.r_State_RNO_1_LC_12_10_4  (
            .in0(N__8562),
            .in1(N__8550),
            .in2(N__8544),
            .in3(N__8541),
            .lcout(),
            .ltout(\Debounce_SW3.r_Count13_0_a7_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_State_LC_12_10_5 .C_ON=1'b0;
    defparam \Debounce_SW3.r_State_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \Debounce_SW3.r_State_LC_12_10_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \Debounce_SW3.r_State_LC_12_10_5  (
            .in0(N__8522),
            .in1(N__8478),
            .in2(N__8502),
            .in3(N__8499),
            .lcout(w_Switch_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8451),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNIOKFA_12_LC_12_10_6 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNIOKFA_12_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNIOKFA_12_LC_12_10_6 .LUT_INIT=16'b0101111101111111;
    LogicCell40 \Debounce_SW3.r_Count_RNIOKFA_12_LC_12_10_6  (
            .in0(N__8299),
            .in1(N__8281),
            .in2(N__8265),
            .in3(N__8245),
            .lcout(),
            .ltout(\Debounce_SW3.un1_r_Count_8lto17_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Debounce_SW3.r_Count_RNI7INF_17_LC_12_10_7 .C_ON=1'b0;
    defparam \Debounce_SW3.r_Count_RNI7INF_17_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \Debounce_SW3.r_Count_RNI7INF_17_LC_12_10_7 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \Debounce_SW3.r_Count_RNI7INF_17_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__8230),
            .in2(N__8217),
            .in3(N__8212),
            .lcout(\Debounce_SW3.un1_r_Count_8lto17_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // State_Machine_Project_Top
